`define STIMULUS_WIDTH      4000
`define DATA_WIDTH			12
`define CTRL_WIDTH			3

module generate_stimuls(y_list, z_list);
    
    output reg [(`DATA_WIDTH * `STIMULUS_WIDTH) - 1 : 0] y_list;
    output reg [(`CTRL_WIDTH * `STIMULUS_WIDTH) - 1 : 0] z_list;

    reg [`DATA_WIDTH - 1 : 0] y[`STIMULUS_WIDTH - 1 : 0];
    reg [`CTRL_WIDTH - 1 : 0] z[`STIMULUS_WIDTH - 1 : 0];

    integer i;

    initial begin
		y[0] = 12'b111001010011;
		z[0] = 3'b110;
		y[1] = 12'b011100010111;
		z[1] = 3'b111;
		y[2] = 12'b000111110001;
		z[2] = 3'b001;
		y[3] = 12'b001000001010;
		z[3] = 3'b011;
		y[4] = 12'b111001110010;
		z[4] = 3'b111;
		y[5] = 12'b000110100010;
		z[5] = 3'b111;
		y[6] = 12'b100111101110;
		z[6] = 3'b011;
		y[7] = 12'b100111101000;
		z[7] = 3'b010;
		y[8] = 12'b010111111001;
		z[8] = 3'b111;
		y[9] = 12'b111101111000;
		z[9] = 3'b111;
		y[10] = 12'b101010011000;
		z[10] = 3'b000;
		y[11] = 12'b011111011101;
		z[11] = 3'b001;
		y[12] = 12'b000101110010;
		z[12] = 3'b110;
		y[13] = 12'b111000001011;
		z[13] = 3'b000;
		y[14] = 12'b111001000001;
		z[14] = 3'b101;
		y[15] = 12'b010100111000;
		z[15] = 3'b000;
		y[16] = 12'b011110110100;
		z[16] = 3'b011;
		y[17] = 12'b110011000001;
		z[17] = 3'b000;
		y[18] = 12'b111100011111;
		z[18] = 3'b000;
		y[19] = 12'b000001100111;
		z[19] = 3'b110;
		y[20] = 12'b000000100101;
		z[20] = 3'b101;
		y[21] = 12'b101011001100;
		z[21] = 3'b001;
		y[22] = 12'b001011101010;
		z[22] = 3'b111;
		y[23] = 12'b101010011011;
		z[23] = 3'b111;
		y[24] = 12'b010010010101;
		z[24] = 3'b110;
		y[25] = 12'b100000101010;
		z[25] = 3'b101;
		y[26] = 12'b101100110001;
		z[26] = 3'b011;
		y[27] = 12'b110001100110;
		z[27] = 3'b101;
		y[28] = 12'b000001001111;
		z[28] = 3'b010;
		y[29] = 12'b101000100100;
		z[29] = 3'b110;
		y[30] = 12'b100110011011;
		z[30] = 3'b010;
		y[31] = 12'b100100101100;
		z[31] = 3'b110;
		y[32] = 12'b110100100001;
		z[32] = 3'b111;
		y[33] = 12'b011111011100;
		z[33] = 3'b111;
		y[34] = 12'b111010000001;
		z[34] = 3'b111;
		y[35] = 12'b100111000000;
		z[35] = 3'b000;
		y[36] = 12'b011101001001;
		z[36] = 3'b100;
		y[37] = 12'b011011100000;
		z[37] = 3'b110;
		y[38] = 12'b101101010110;
		z[38] = 3'b111;
		y[39] = 12'b101110000011;
		z[39] = 3'b011;
		y[40] = 12'b000110001111;
		z[40] = 3'b111;
		y[41] = 12'b001011010110;
		z[41] = 3'b100;
		y[42] = 12'b111111111110;
		z[42] = 3'b000;
		y[43] = 12'b100000011100;
		z[43] = 3'b100;
		y[44] = 12'b010111001110;
		z[44] = 3'b011;
		y[45] = 12'b010100100010;
		z[45] = 3'b101;
		y[46] = 12'b100101001011;
		z[46] = 3'b011;
		y[47] = 12'b100010010011;
		z[47] = 3'b100;
		y[48] = 12'b001001110111;
		z[48] = 3'b011;
		y[49] = 12'b111010100101;
		z[49] = 3'b110;
		y[50] = 12'b001110110101;
		z[50] = 3'b101;
		y[51] = 12'b111111011100;
		z[51] = 3'b000;
		y[52] = 12'b101100001011;
		z[52] = 3'b110;
		y[53] = 12'b111010110111;
		z[53] = 3'b111;
		y[54] = 12'b100111111100;
		z[54] = 3'b000;
		y[55] = 12'b110010000010;
		z[55] = 3'b000;
		y[56] = 12'b110010100100;
		z[56] = 3'b111;
		y[57] = 12'b001000011100;
		z[57] = 3'b110;
		y[58] = 12'b110101111000;
		z[58] = 3'b001;
		y[59] = 12'b100010000001;
		z[59] = 3'b110;
		y[60] = 12'b011000111011;
		z[60] = 3'b001;
		y[61] = 12'b111101011010;
		z[61] = 3'b000;
		y[62] = 12'b000110011000;
		z[62] = 3'b000;
		y[63] = 12'b000011010100;
		z[63] = 3'b101;
		y[64] = 12'b011001001101;
		z[64] = 3'b100;
		y[65] = 12'b000100000100;
		z[65] = 3'b100;
		y[66] = 12'b000110001110;
		z[66] = 3'b011;
		y[67] = 12'b111101000110;
		z[67] = 3'b101;
		y[68] = 12'b000010000010;
		z[68] = 3'b101;
		y[69] = 12'b101111011001;
		z[69] = 3'b011;
		y[70] = 12'b001011011001;
		z[70] = 3'b001;
		y[71] = 12'b010110000010;
		z[71] = 3'b110;
		y[72] = 12'b010000001111;
		z[72] = 3'b000;
		y[73] = 12'b101111011001;
		z[73] = 3'b100;
		y[74] = 12'b100111111010;
		z[74] = 3'b101;
		y[75] = 12'b011100010111;
		z[75] = 3'b000;
		y[76] = 12'b100111010100;
		z[76] = 3'b000;
		y[77] = 12'b010001001000;
		z[77] = 3'b011;
		y[78] = 12'b001100000101;
		z[78] = 3'b001;
		y[79] = 12'b011101001001;
		z[79] = 3'b111;
		y[80] = 12'b100001001011;
		z[80] = 3'b000;
		y[81] = 12'b110101000010;
		z[81] = 3'b101;
		y[82] = 12'b000011100101;
		z[82] = 3'b011;
		y[83] = 12'b011101000110;
		z[83] = 3'b000;
		y[84] = 12'b100000111111;
		z[84] = 3'b011;
		y[85] = 12'b001010011010;
		z[85] = 3'b000;
		y[86] = 12'b100111001011;
		z[86] = 3'b001;
		y[87] = 12'b001010110100;
		z[87] = 3'b100;
		y[88] = 12'b100110011101;
		z[88] = 3'b011;
		y[89] = 12'b000000100000;
		z[89] = 3'b000;
		y[90] = 12'b111111000011;
		z[90] = 3'b001;
		y[91] = 12'b111111001011;
		z[91] = 3'b000;
		y[92] = 12'b010000111011;
		z[92] = 3'b011;
		y[93] = 12'b101000001111;
		z[93] = 3'b001;
		y[94] = 12'b100111010010;
		z[94] = 3'b001;
		y[95] = 12'b111010011000;
		z[95] = 3'b101;
		y[96] = 12'b000110100110;
		z[96] = 3'b111;
		y[97] = 12'b000011111100;
		z[97] = 3'b011;
		y[98] = 12'b110000010001;
		z[98] = 3'b101;
		y[99] = 12'b100110000000;
		z[99] = 3'b010;
		y[100] = 12'b111011110000;
		z[100] = 3'b110;
		y[101] = 12'b001110100101;
		z[101] = 3'b110;
		y[102] = 12'b010110110110;
		z[102] = 3'b011;
		y[103] = 12'b111000000001;
		z[103] = 3'b110;
		y[104] = 12'b000010010110;
		z[104] = 3'b001;
		y[105] = 12'b011010010101;
		z[105] = 3'b011;
		y[106] = 12'b110001001101;
		z[106] = 3'b010;
		y[107] = 12'b000110010000;
		z[107] = 3'b011;
		y[108] = 12'b100101100111;
		z[108] = 3'b100;
		y[109] = 12'b110010000001;
		z[109] = 3'b000;
		y[110] = 12'b101110010011;
		z[110] = 3'b110;
		y[111] = 12'b101010110111;
		z[111] = 3'b110;
		y[112] = 12'b111000101001;
		z[112] = 3'b010;
		y[113] = 12'b010011000011;
		z[113] = 3'b101;
		y[114] = 12'b000111010111;
		z[114] = 3'b111;
		y[115] = 12'b101110011000;
		z[115] = 3'b101;
		y[116] = 12'b111100001110;
		z[116] = 3'b101;
		y[117] = 12'b010010110000;
		z[117] = 3'b001;
		y[118] = 12'b111000010001;
		z[118] = 3'b100;
		y[119] = 12'b001011111001;
		z[119] = 3'b010;
		y[120] = 12'b010010101101;
		z[120] = 3'b110;
		y[121] = 12'b100010100000;
		z[121] = 3'b000;
		y[122] = 12'b010111011101;
		z[122] = 3'b010;
		y[123] = 12'b111001001010;
		z[123] = 3'b100;
		y[124] = 12'b001011100100;
		z[124] = 3'b110;
		y[125] = 12'b100001100000;
		z[125] = 3'b010;
		y[126] = 12'b010000111010;
		z[126] = 3'b110;
		y[127] = 12'b100001010000;
		z[127] = 3'b100;
		y[128] = 12'b100101101001;
		z[128] = 3'b110;
		y[129] = 12'b100010111100;
		z[129] = 3'b011;
		y[130] = 12'b111100010010;
		z[130] = 3'b000;
		y[131] = 12'b001110010000;
		z[131] = 3'b011;
		y[132] = 12'b000010011011;
		z[132] = 3'b011;
		y[133] = 12'b101000111011;
		z[133] = 3'b011;
		y[134] = 12'b111010101000;
		z[134] = 3'b100;
		y[135] = 12'b110001100010;
		z[135] = 3'b011;
		y[136] = 12'b010010000111;
		z[136] = 3'b011;
		y[137] = 12'b110011101010;
		z[137] = 3'b001;
		y[138] = 12'b111111001111;
		z[138] = 3'b101;
		y[139] = 12'b011110111100;
		z[139] = 3'b100;
		y[140] = 12'b101000001111;
		z[140] = 3'b010;
		y[141] = 12'b101110011000;
		z[141] = 3'b001;
		y[142] = 12'b110111101101;
		z[142] = 3'b111;
		y[143] = 12'b011011110111;
		z[143] = 3'b101;
		y[144] = 12'b110101111011;
		z[144] = 3'b001;
		y[145] = 12'b110000000110;
		z[145] = 3'b000;
		y[146] = 12'b110111101111;
		z[146] = 3'b101;
		y[147] = 12'b101110010111;
		z[147] = 3'b001;
		y[148] = 12'b011111010101;
		z[148] = 3'b000;
		y[149] = 12'b001000001111;
		z[149] = 3'b100;
		y[150] = 12'b111011100000;
		z[150] = 3'b000;
		y[151] = 12'b010110000000;
		z[151] = 3'b011;
		y[152] = 12'b110110000011;
		z[152] = 3'b111;
		y[153] = 12'b001011101101;
		z[153] = 3'b111;
		y[154] = 12'b110101111001;
		z[154] = 3'b100;
		y[155] = 12'b101011010001;
		z[155] = 3'b001;
		y[156] = 12'b101001101011;
		z[156] = 3'b011;
		y[157] = 12'b101011100101;
		z[157] = 3'b111;
		y[158] = 12'b010001101001;
		z[158] = 3'b111;
		y[159] = 12'b010101000011;
		z[159] = 3'b000;
		y[160] = 12'b100010011110;
		z[160] = 3'b001;
		y[161] = 12'b100000011111;
		z[161] = 3'b011;
		y[162] = 12'b010010000100;
		z[162] = 3'b100;
		y[163] = 12'b010111010011;
		z[163] = 3'b100;
		y[164] = 12'b101100111110;
		z[164] = 3'b100;
		y[165] = 12'b111000100100;
		z[165] = 3'b011;
		y[166] = 12'b100011001101;
		z[166] = 3'b110;
		y[167] = 12'b100111110101;
		z[167] = 3'b110;
		y[168] = 12'b001010111001;
		z[168] = 3'b100;
		y[169] = 12'b000110110000;
		z[169] = 3'b001;
		y[170] = 12'b001101111110;
		z[170] = 3'b100;
		y[171] = 12'b000101111010;
		z[171] = 3'b101;
		y[172] = 12'b100100100000;
		z[172] = 3'b011;
		y[173] = 12'b011100101000;
		z[173] = 3'b001;
		y[174] = 12'b000010111110;
		z[174] = 3'b011;
		y[175] = 12'b111000110000;
		z[175] = 3'b100;
		y[176] = 12'b111011100001;
		z[176] = 3'b000;
		y[177] = 12'b110111010010;
		z[177] = 3'b010;
		y[178] = 12'b011001011011;
		z[178] = 3'b010;
		y[179] = 12'b010111000111;
		z[179] = 3'b001;
		y[180] = 12'b111110100101;
		z[180] = 3'b010;
		y[181] = 12'b001100111100;
		z[181] = 3'b000;
		y[182] = 12'b010001100011;
		z[182] = 3'b110;
		y[183] = 12'b100001100000;
		z[183] = 3'b100;
		y[184] = 12'b110110100000;
		z[184] = 3'b001;
		y[185] = 12'b000100100001;
		z[185] = 3'b101;
		y[186] = 12'b001110001010;
		z[186] = 3'b100;
		y[187] = 12'b000111011100;
		z[187] = 3'b101;
		y[188] = 12'b010110100010;
		z[188] = 3'b110;
		y[189] = 12'b000010000111;
		z[189] = 3'b000;
		y[190] = 12'b000111010011;
		z[190] = 3'b010;
		y[191] = 12'b010100000000;
		z[191] = 3'b010;
		y[192] = 12'b110100100001;
		z[192] = 3'b110;
		y[193] = 12'b101000010001;
		z[193] = 3'b111;
		y[194] = 12'b111000011111;
		z[194] = 3'b011;
		y[195] = 12'b100000101010;
		z[195] = 3'b101;
		y[196] = 12'b010100001000;
		z[196] = 3'b001;
		y[197] = 12'b010010101001;
		z[197] = 3'b000;
		y[198] = 12'b001000101110;
		z[198] = 3'b001;
		y[199] = 12'b101001101101;
		z[199] = 3'b110;
		y[200] = 12'b011100011110;
		z[200] = 3'b111;
		y[201] = 12'b100001101100;
		z[201] = 3'b100;
		y[202] = 12'b001101000010;
		z[202] = 3'b111;
		y[203] = 12'b100000110001;
		z[203] = 3'b000;
		y[204] = 12'b111010111001;
		z[204] = 3'b101;
		y[205] = 12'b011010011001;
		z[205] = 3'b101;
		y[206] = 12'b100000111100;
		z[206] = 3'b011;
		y[207] = 12'b001010011000;
		z[207] = 3'b010;
		y[208] = 12'b010100010111;
		z[208] = 3'b000;
		y[209] = 12'b010100110100;
		z[209] = 3'b001;
		y[210] = 12'b010100010101;
		z[210] = 3'b111;
		y[211] = 12'b101001110110;
		z[211] = 3'b110;
		y[212] = 12'b010100010101;
		z[212] = 3'b110;
		y[213] = 12'b100001110000;
		z[213] = 3'b101;
		y[214] = 12'b100000111101;
		z[214] = 3'b101;
		y[215] = 12'b101001100110;
		z[215] = 3'b011;
		y[216] = 12'b110000001001;
		z[216] = 3'b110;
		y[217] = 12'b100101101110;
		z[217] = 3'b110;
		y[218] = 12'b100010010011;
		z[218] = 3'b100;
		y[219] = 12'b000101001011;
		z[219] = 3'b110;
		y[220] = 12'b000010000010;
		z[220] = 3'b101;
		y[221] = 12'b000100000100;
		z[221] = 3'b100;
		y[222] = 12'b100001111000;
		z[222] = 3'b110;
		y[223] = 12'b001111011100;
		z[223] = 3'b101;
		y[224] = 12'b100100110000;
		z[224] = 3'b100;
		y[225] = 12'b100001100010;
		z[225] = 3'b001;
		y[226] = 12'b100011011100;
		z[226] = 3'b110;
		y[227] = 12'b011100100100;
		z[227] = 3'b101;
		y[228] = 12'b100001001100;
		z[228] = 3'b010;
		y[229] = 12'b010101101111;
		z[229] = 3'b010;
		y[230] = 12'b000011111111;
		z[230] = 3'b111;
		y[231] = 12'b101010100101;
		z[231] = 3'b011;
		y[232] = 12'b011000100010;
		z[232] = 3'b011;
		y[233] = 12'b000001001100;
		z[233] = 3'b010;
		y[234] = 12'b110110011111;
		z[234] = 3'b111;
		y[235] = 12'b011000110111;
		z[235] = 3'b100;
		y[236] = 12'b110111111011;
		z[236] = 3'b100;
		y[237] = 12'b101100001100;
		z[237] = 3'b000;
		y[238] = 12'b110000111001;
		z[238] = 3'b011;
		y[239] = 12'b101000010110;
		z[239] = 3'b110;
		y[240] = 12'b011110111010;
		z[240] = 3'b000;
		y[241] = 12'b110010100000;
		z[241] = 3'b001;
		y[242] = 12'b110000101011;
		z[242] = 3'b100;
		y[243] = 12'b010001001011;
		z[243] = 3'b100;
		y[244] = 12'b010011011110;
		z[244] = 3'b011;
		y[245] = 12'b101010111100;
		z[245] = 3'b100;
		y[246] = 12'b101000011010;
		z[246] = 3'b000;
		y[247] = 12'b110001000100;
		z[247] = 3'b101;
		y[248] = 12'b011110110000;
		z[248] = 3'b110;
		y[249] = 12'b000001010111;
		z[249] = 3'b000;
		y[250] = 12'b101111110100;
		z[250] = 3'b000;
		y[251] = 12'b011110110000;
		z[251] = 3'b101;
		y[252] = 12'b110011011100;
		z[252] = 3'b100;
		y[253] = 12'b000010000101;
		z[253] = 3'b110;
		y[254] = 12'b010110110101;
		z[254] = 3'b001;
		y[255] = 12'b101001110111;
		z[255] = 3'b001;
		y[256] = 12'b100101100100;
		z[256] = 3'b110;
		y[257] = 12'b001011011111;
		z[257] = 3'b000;
		y[258] = 12'b100010011101;
		z[258] = 3'b001;
		y[259] = 12'b111111110001;
		z[259] = 3'b010;
		y[260] = 12'b011010110110;
		z[260] = 3'b000;
		y[261] = 12'b011001100111;
		z[261] = 3'b001;
		y[262] = 12'b100000010101;
		z[262] = 3'b011;
		y[263] = 12'b110100100110;
		z[263] = 3'b111;
		y[264] = 12'b111000001000;
		z[264] = 3'b100;
		y[265] = 12'b000010100011;
		z[265] = 3'b011;
		y[266] = 12'b101001100110;
		z[266] = 3'b001;
		y[267] = 12'b000111001111;
		z[267] = 3'b100;
		y[268] = 12'b001101000111;
		z[268] = 3'b010;
		y[269] = 12'b101011000001;
		z[269] = 3'b100;
		y[270] = 12'b111100100011;
		z[270] = 3'b000;
		y[271] = 12'b000111110010;
		z[271] = 3'b001;
		y[272] = 12'b100001011111;
		z[272] = 3'b011;
		y[273] = 12'b100101111100;
		z[273] = 3'b101;
		y[274] = 12'b110110011011;
		z[274] = 3'b111;
		y[275] = 12'b001010110111;
		z[275] = 3'b111;
		y[276] = 12'b011100101101;
		z[276] = 3'b000;
		y[277] = 12'b101101000000;
		z[277] = 3'b000;
		y[278] = 12'b100011011000;
		z[278] = 3'b110;
		y[279] = 12'b010000010000;
		z[279] = 3'b011;
		y[280] = 12'b101001110101;
		z[280] = 3'b000;
		y[281] = 12'b111110111001;
		z[281] = 3'b011;
		y[282] = 12'b111110111000;
		z[282] = 3'b111;
		y[283] = 12'b001111110010;
		z[283] = 3'b010;
		y[284] = 12'b000100001101;
		z[284] = 3'b000;
		y[285] = 12'b111011011011;
		z[285] = 3'b111;
		y[286] = 12'b010101101000;
		z[286] = 3'b111;
		y[287] = 12'b100000001101;
		z[287] = 3'b110;
		y[288] = 12'b000101001000;
		z[288] = 3'b110;
		y[289] = 12'b011100011100;
		z[289] = 3'b011;
		y[290] = 12'b010001011011;
		z[290] = 3'b001;
		y[291] = 12'b011110010000;
		z[291] = 3'b110;
		y[292] = 12'b110000110111;
		z[292] = 3'b110;
		y[293] = 12'b011001110111;
		z[293] = 3'b110;
		y[294] = 12'b010000001110;
		z[294] = 3'b100;
		y[295] = 12'b100001101000;
		z[295] = 3'b101;
		y[296] = 12'b111010101011;
		z[296] = 3'b000;
		y[297] = 12'b011110000011;
		z[297] = 3'b111;
		y[298] = 12'b101011000101;
		z[298] = 3'b110;
		y[299] = 12'b010001100001;
		z[299] = 3'b011;
		y[300] = 12'b011110001010;
		z[300] = 3'b101;
		y[301] = 12'b111000110110;
		z[301] = 3'b000;
		y[302] = 12'b101010011100;
		z[302] = 3'b001;
		y[303] = 12'b111100001110;
		z[303] = 3'b000;
		y[304] = 12'b011001001111;
		z[304] = 3'b111;
		y[305] = 12'b001100110000;
		z[305] = 3'b001;
		y[306] = 12'b111001111110;
		z[306] = 3'b001;
		y[307] = 12'b010000010111;
		z[307] = 3'b110;
		y[308] = 12'b110101110111;
		z[308] = 3'b010;
		y[309] = 12'b100110011010;
		z[309] = 3'b010;
		y[310] = 12'b111010000010;
		z[310] = 3'b000;
		y[311] = 12'b011011001000;
		z[311] = 3'b000;
		y[312] = 12'b000010001001;
		z[312] = 3'b101;
		y[313] = 12'b110001000111;
		z[313] = 3'b110;
		y[314] = 12'b000011101010;
		z[314] = 3'b110;
		y[315] = 12'b000100011111;
		z[315] = 3'b100;
		y[316] = 12'b011001011010;
		z[316] = 3'b110;
		y[317] = 12'b101010110110;
		z[317] = 3'b011;
		y[318] = 12'b010000011000;
		z[318] = 3'b011;
		y[319] = 12'b011010010100;
		z[319] = 3'b010;
		y[320] = 12'b100010110111;
		z[320] = 3'b001;
		y[321] = 12'b011101001100;
		z[321] = 3'b001;
		y[322] = 12'b010110000001;
		z[322] = 3'b000;
		y[323] = 12'b100010101111;
		z[323] = 3'b110;
		y[324] = 12'b110000111110;
		z[324] = 3'b111;
		y[325] = 12'b101110111111;
		z[325] = 3'b010;
		y[326] = 12'b100100110100;
		z[326] = 3'b110;
		y[327] = 12'b111001011001;
		z[327] = 3'b000;
		y[328] = 12'b011100101010;
		z[328] = 3'b001;
		y[329] = 12'b101010011001;
		z[329] = 3'b011;
		y[330] = 12'b001010001001;
		z[330] = 3'b000;
		y[331] = 12'b111001111000;
		z[331] = 3'b111;
		y[332] = 12'b011100100111;
		z[332] = 3'b011;
		y[333] = 12'b000000110100;
		z[333] = 3'b111;
		y[334] = 12'b001010101101;
		z[334] = 3'b011;
		y[335] = 12'b011100010010;
		z[335] = 3'b100;
		y[336] = 12'b000111010111;
		z[336] = 3'b111;
		y[337] = 12'b100110011000;
		z[337] = 3'b010;
		y[338] = 12'b111111001101;
		z[338] = 3'b111;
		y[339] = 12'b000101001111;
		z[339] = 3'b111;
		y[340] = 12'b101101101011;
		z[340] = 3'b001;
		y[341] = 12'b000111101001;
		z[341] = 3'b011;
		y[342] = 12'b100100010110;
		z[342] = 3'b111;
		y[343] = 12'b100011011100;
		z[343] = 3'b100;
		y[344] = 12'b110110011011;
		z[344] = 3'b011;
		y[345] = 12'b101000111011;
		z[345] = 3'b101;
		y[346] = 12'b011110000001;
		z[346] = 3'b000;
		y[347] = 12'b101101100100;
		z[347] = 3'b011;
		y[348] = 12'b010101111101;
		z[348] = 3'b111;
		y[349] = 12'b111100001001;
		z[349] = 3'b000;
		y[350] = 12'b101000000110;
		z[350] = 3'b111;
		y[351] = 12'b000101111001;
		z[351] = 3'b011;
		y[352] = 12'b000011110010;
		z[352] = 3'b000;
		y[353] = 12'b101010110000;
		z[353] = 3'b010;
		y[354] = 12'b001001101100;
		z[354] = 3'b010;
		y[355] = 12'b010100011110;
		z[355] = 3'b110;
		y[356] = 12'b000000101011;
		z[356] = 3'b101;
		y[357] = 12'b000000101101;
		z[357] = 3'b001;
		y[358] = 12'b100111100001;
		z[358] = 3'b111;
		y[359] = 12'b100111101110;
		z[359] = 3'b010;
		y[360] = 12'b100110110001;
		z[360] = 3'b111;
		y[361] = 12'b010110110101;
		z[361] = 3'b001;
		y[362] = 12'b101111001010;
		z[362] = 3'b100;
		y[363] = 12'b101010101101;
		z[363] = 3'b011;
		y[364] = 12'b101101110000;
		z[364] = 3'b011;
		y[365] = 12'b000001010111;
		z[365] = 3'b011;
		y[366] = 12'b000010011111;
		z[366] = 3'b110;
		y[367] = 12'b011111010001;
		z[367] = 3'b001;
		y[368] = 12'b011111101001;
		z[368] = 3'b001;
		y[369] = 12'b001111010110;
		z[369] = 3'b001;
		y[370] = 12'b110100100100;
		z[370] = 3'b101;
		y[371] = 12'b010010010100;
		z[371] = 3'b001;
		y[372] = 12'b101011110100;
		z[372] = 3'b011;
		y[373] = 12'b111100101100;
		z[373] = 3'b001;
		y[374] = 12'b001010111111;
		z[374] = 3'b110;
		y[375] = 12'b111100110001;
		z[375] = 3'b111;
		y[376] = 12'b001100001111;
		z[376] = 3'b010;
		y[377] = 12'b110001101010;
		z[377] = 3'b110;
		y[378] = 12'b110011000011;
		z[378] = 3'b101;
		y[379] = 12'b000111101100;
		z[379] = 3'b111;
		y[380] = 12'b110100011101;
		z[380] = 3'b111;
		y[381] = 12'b001010110110;
		z[381] = 3'b010;
		y[382] = 12'b010010101011;
		z[382] = 3'b011;
		y[383] = 12'b000001111010;
		z[383] = 3'b100;
		y[384] = 12'b101010010001;
		z[384] = 3'b111;
		y[385] = 12'b011011011111;
		z[385] = 3'b110;
		y[386] = 12'b101011000110;
		z[386] = 3'b110;
		y[387] = 12'b011000011110;
		z[387] = 3'b110;
		y[388] = 12'b101100110101;
		z[388] = 3'b100;
		y[389] = 12'b001110000001;
		z[389] = 3'b111;
		y[390] = 12'b010011101010;
		z[390] = 3'b101;
		y[391] = 12'b011011101000;
		z[391] = 3'b000;
		y[392] = 12'b110011011001;
		z[392] = 3'b011;
		y[393] = 12'b010000001001;
		z[393] = 3'b111;
		y[394] = 12'b110111100110;
		z[394] = 3'b101;
		y[395] = 12'b001100010000;
		z[395] = 3'b101;
		y[396] = 12'b111011000100;
		z[396] = 3'b010;
		y[397] = 12'b000011110111;
		z[397] = 3'b000;
		y[398] = 12'b101101101101;
		z[398] = 3'b111;
		y[399] = 12'b111101100100;
		z[399] = 3'b001;
		y[400] = 12'b100110111110;
		z[400] = 3'b000;
		y[401] = 12'b100001111110;
		z[401] = 3'b000;
		y[402] = 12'b111010100000;
		z[402] = 3'b110;
		y[403] = 12'b000011010100;
		z[403] = 3'b100;
		y[404] = 12'b100011101000;
		z[404] = 3'b101;
		y[405] = 12'b010101101110;
		z[405] = 3'b110;
		y[406] = 12'b111010101101;
		z[406] = 3'b110;
		y[407] = 12'b111101100110;
		z[407] = 3'b011;
		y[408] = 12'b001001011001;
		z[408] = 3'b010;
		y[409] = 12'b100110000111;
		z[409] = 3'b101;
		y[410] = 12'b011001111010;
		z[410] = 3'b110;
		y[411] = 12'b011110101111;
		z[411] = 3'b000;
		y[412] = 12'b110110100110;
		z[412] = 3'b010;
		y[413] = 12'b011000011000;
		z[413] = 3'b000;
		y[414] = 12'b011101011011;
		z[414] = 3'b010;
		y[415] = 12'b100010010100;
		z[415] = 3'b110;
		y[416] = 12'b111100000111;
		z[416] = 3'b100;
		y[417] = 12'b100011001011;
		z[417] = 3'b000;
		y[418] = 12'b100110111100;
		z[418] = 3'b011;
		y[419] = 12'b001000111010;
		z[419] = 3'b000;
		y[420] = 12'b001100000010;
		z[420] = 3'b011;
		y[421] = 12'b111111001100;
		z[421] = 3'b010;
		y[422] = 12'b011011001011;
		z[422] = 3'b011;
		y[423] = 12'b111010111111;
		z[423] = 3'b100;
		y[424] = 12'b110110100011;
		z[424] = 3'b011;
		y[425] = 12'b011101101001;
		z[425] = 3'b110;
		y[426] = 12'b001011101101;
		z[426] = 3'b111;
		y[427] = 12'b101000110010;
		z[427] = 3'b111;
		y[428] = 12'b010001010100;
		z[428] = 3'b010;
		y[429] = 12'b001001110000;
		z[429] = 3'b001;
		y[430] = 12'b110011111111;
		z[430] = 3'b001;
		y[431] = 12'b101101000100;
		z[431] = 3'b110;
		y[432] = 12'b001001101111;
		z[432] = 3'b110;
		y[433] = 12'b011110010010;
		z[433] = 3'b010;
		y[434] = 12'b101010111001;
		z[434] = 3'b010;
		y[435] = 12'b110111100110;
		z[435] = 3'b010;
		y[436] = 12'b100110110100;
		z[436] = 3'b001;
		y[437] = 12'b101110001100;
		z[437] = 3'b111;
		y[438] = 12'b011100000100;
		z[438] = 3'b011;
		y[439] = 12'b100011010001;
		z[439] = 3'b111;
		y[440] = 12'b001010100010;
		z[440] = 3'b110;
		y[441] = 12'b000001100100;
		z[441] = 3'b010;
		y[442] = 12'b001110010010;
		z[442] = 3'b011;
		y[443] = 12'b100101101100;
		z[443] = 3'b110;
		y[444] = 12'b011101110101;
		z[444] = 3'b111;
		y[445] = 12'b010000010111;
		z[445] = 3'b100;
		y[446] = 12'b101000000111;
		z[446] = 3'b011;
		y[447] = 12'b101100101101;
		z[447] = 3'b110;
		y[448] = 12'b010000000101;
		z[448] = 3'b011;
		y[449] = 12'b001010010011;
		z[449] = 3'b111;
		y[450] = 12'b011110011110;
		z[450] = 3'b001;
		y[451] = 12'b001111011100;
		z[451] = 3'b000;
		y[452] = 12'b000110010001;
		z[452] = 3'b001;
		y[453] = 12'b011100001001;
		z[453] = 3'b000;
		y[454] = 12'b100111101010;
		z[454] = 3'b100;
		y[455] = 12'b000000111010;
		z[455] = 3'b010;
		y[456] = 12'b000000111100;
		z[456] = 3'b000;
		y[457] = 12'b011111110111;
		z[457] = 3'b100;
		y[458] = 12'b001011010010;
		z[458] = 3'b100;
		y[459] = 12'b110100111011;
		z[459] = 3'b010;
		y[460] = 12'b010000001000;
		z[460] = 3'b001;
		y[461] = 12'b000011110010;
		z[461] = 3'b101;
		y[462] = 12'b110101111000;
		z[462] = 3'b010;
		y[463] = 12'b101110000010;
		z[463] = 3'b010;
		y[464] = 12'b000010010000;
		z[464] = 3'b101;
		y[465] = 12'b111010011001;
		z[465] = 3'b011;
		y[466] = 12'b010001000100;
		z[466] = 3'b000;
		y[467] = 12'b000100011000;
		z[467] = 3'b110;
		y[468] = 12'b110110110000;
		z[468] = 3'b011;
		y[469] = 12'b000000101011;
		z[469] = 3'b001;
		y[470] = 12'b100100110110;
		z[470] = 3'b111;
		y[471] = 12'b101111101010;
		z[471] = 3'b101;
		y[472] = 12'b101011100001;
		z[472] = 3'b100;
		y[473] = 12'b010101110111;
		z[473] = 3'b001;
		y[474] = 12'b001100111101;
		z[474] = 3'b111;
		y[475] = 12'b111010101100;
		z[475] = 3'b000;
		y[476] = 12'b011110100001;
		z[476] = 3'b101;
		y[477] = 12'b001110110111;
		z[477] = 3'b001;
		y[478] = 12'b101100110100;
		z[478] = 3'b111;
		y[479] = 12'b011010110001;
		z[479] = 3'b100;
		y[480] = 12'b011100110000;
		z[480] = 3'b011;
		y[481] = 12'b110001011010;
		z[481] = 3'b100;
		y[482] = 12'b001111111110;
		z[482] = 3'b110;
		y[483] = 12'b101101111010;
		z[483] = 3'b011;
		y[484] = 12'b101100000100;
		z[484] = 3'b100;
		y[485] = 12'b001001111111;
		z[485] = 3'b000;
		y[486] = 12'b010000010011;
		z[486] = 3'b011;
		y[487] = 12'b011011100001;
		z[487] = 3'b111;
		y[488] = 12'b101001110010;
		z[488] = 3'b101;
		y[489] = 12'b011100000010;
		z[489] = 3'b110;
		y[490] = 12'b111010110110;
		z[490] = 3'b011;
		y[491] = 12'b100100011110;
		z[491] = 3'b110;
		y[492] = 12'b010010010101;
		z[492] = 3'b010;
		y[493] = 12'b100011101111;
		z[493] = 3'b011;
		y[494] = 12'b001110011000;
		z[494] = 3'b111;
		y[495] = 12'b111001000101;
		z[495] = 3'b110;
		y[496] = 12'b001001011011;
		z[496] = 3'b101;
		y[497] = 12'b111100000110;
		z[497] = 3'b100;
		y[498] = 12'b110000001000;
		z[498] = 3'b000;
		y[499] = 12'b000001000100;
		z[499] = 3'b101;
		y[500] = 12'b111100010111;
		z[500] = 3'b110;
		y[501] = 12'b101110001000;
		z[501] = 3'b101;
		y[502] = 12'b001010000000;
		z[502] = 3'b001;
		y[503] = 12'b110101001100;
		z[503] = 3'b010;
		y[504] = 12'b101011111000;
		z[504] = 3'b011;
		y[505] = 12'b011011001110;
		z[505] = 3'b101;
		y[506] = 12'b110000001000;
		z[506] = 3'b110;
		y[507] = 12'b001011111100;
		z[507] = 3'b010;
		y[508] = 12'b010010111010;
		z[508] = 3'b100;
		y[509] = 12'b001101111010;
		z[509] = 3'b000;
		y[510] = 12'b110100111111;
		z[510] = 3'b111;
		y[511] = 12'b101010111110;
		z[511] = 3'b101;
		y[512] = 12'b111000100001;
		z[512] = 3'b011;
		y[513] = 12'b010100111100;
		z[513] = 3'b000;
		y[514] = 12'b001100111001;
		z[514] = 3'b001;
		y[515] = 12'b010000111000;
		z[515] = 3'b011;
		y[516] = 12'b101110111100;
		z[516] = 3'b110;
		y[517] = 12'b011110011100;
		z[517] = 3'b001;
		y[518] = 12'b111101001010;
		z[518] = 3'b110;
		y[519] = 12'b010011111111;
		z[519] = 3'b100;
		y[520] = 12'b101001111110;
		z[520] = 3'b101;
		y[521] = 12'b101010011001;
		z[521] = 3'b000;
		y[522] = 12'b101001001000;
		z[522] = 3'b110;
		y[523] = 12'b000101010111;
		z[523] = 3'b101;
		y[524] = 12'b101100100001;
		z[524] = 3'b110;
		y[525] = 12'b010111011010;
		z[525] = 3'b011;
		y[526] = 12'b010000011001;
		z[526] = 3'b010;
		y[527] = 12'b100110111101;
		z[527] = 3'b011;
		y[528] = 12'b110011111101;
		z[528] = 3'b101;
		y[529] = 12'b101111001001;
		z[529] = 3'b000;
		y[530] = 12'b001110100110;
		z[530] = 3'b011;
		y[531] = 12'b010110111110;
		z[531] = 3'b101;
		y[532] = 12'b001011101110;
		z[532] = 3'b111;
		y[533] = 12'b111010011000;
		z[533] = 3'b110;
		y[534] = 12'b000101101011;
		z[534] = 3'b110;
		y[535] = 12'b000111101000;
		z[535] = 3'b100;
		y[536] = 12'b100100110011;
		z[536] = 3'b111;
		y[537] = 12'b100110110100;
		z[537] = 3'b101;
		y[538] = 12'b010000101010;
		z[538] = 3'b000;
		y[539] = 12'b000111100110;
		z[539] = 3'b100;
		y[540] = 12'b000011111000;
		z[540] = 3'b100;
		y[541] = 12'b101010101110;
		z[541] = 3'b110;
		y[542] = 12'b000000111011;
		z[542] = 3'b111;
		y[543] = 12'b011011011001;
		z[543] = 3'b001;
		y[544] = 12'b111111010110;
		z[544] = 3'b100;
		y[545] = 12'b010001011100;
		z[545] = 3'b101;
		y[546] = 12'b101010101000;
		z[546] = 3'b110;
		y[547] = 12'b111110111100;
		z[547] = 3'b000;
		y[548] = 12'b100011110101;
		z[548] = 3'b101;
		y[549] = 12'b010101101110;
		z[549] = 3'b100;
		y[550] = 12'b100111000101;
		z[550] = 3'b010;
		y[551] = 12'b001110001110;
		z[551] = 3'b000;
		y[552] = 12'b101010000011;
		z[552] = 3'b010;
		y[553] = 12'b000010101001;
		z[553] = 3'b110;
		y[554] = 12'b110011010101;
		z[554] = 3'b000;
		y[555] = 12'b000110001100;
		z[555] = 3'b001;
		y[556] = 12'b010100000001;
		z[556] = 3'b010;
		y[557] = 12'b010010011100;
		z[557] = 3'b110;
		y[558] = 12'b100010111100;
		z[558] = 3'b111;
		y[559] = 12'b100001011110;
		z[559] = 3'b010;
		y[560] = 12'b000000100010;
		z[560] = 3'b101;
		y[561] = 12'b000000000110;
		z[561] = 3'b111;
		y[562] = 12'b011000111101;
		z[562] = 3'b101;
		y[563] = 12'b111001100001;
		z[563] = 3'b111;
		y[564] = 12'b011000010001;
		z[564] = 3'b111;
		y[565] = 12'b111101001100;
		z[565] = 3'b100;
		y[566] = 12'b010110101100;
		z[566] = 3'b001;
		y[567] = 12'b110110111010;
		z[567] = 3'b011;
		y[568] = 12'b110001101010;
		z[568] = 3'b101;
		y[569] = 12'b011100100001;
		z[569] = 3'b000;
		y[570] = 12'b011011101111;
		z[570] = 3'b001;
		y[571] = 12'b011101101100;
		z[571] = 3'b011;
		y[572] = 12'b100100111111;
		z[572] = 3'b011;
		y[573] = 12'b001011001010;
		z[573] = 3'b100;
		y[574] = 12'b100101001101;
		z[574] = 3'b001;
		y[575] = 12'b101111110101;
		z[575] = 3'b110;
		y[576] = 12'b110000000110;
		z[576] = 3'b010;
		y[577] = 12'b111101010000;
		z[577] = 3'b011;
		y[578] = 12'b000001101111;
		z[578] = 3'b110;
		y[579] = 12'b011010001000;
		z[579] = 3'b101;
		y[580] = 12'b111101110000;
		z[580] = 3'b000;
		y[581] = 12'b101100000011;
		z[581] = 3'b011;
		y[582] = 12'b101000011011;
		z[582] = 3'b001;
		y[583] = 12'b100101101000;
		z[583] = 3'b111;
		y[584] = 12'b010101000011;
		z[584] = 3'b011;
		y[585] = 12'b100110111000;
		z[585] = 3'b101;
		y[586] = 12'b001000011111;
		z[586] = 3'b011;
		y[587] = 12'b100010111111;
		z[587] = 3'b000;
		y[588] = 12'b001100111001;
		z[588] = 3'b111;
		y[589] = 12'b111010011001;
		z[589] = 3'b110;
		y[590] = 12'b011111010101;
		z[590] = 3'b100;
		y[591] = 12'b001100110010;
		z[591] = 3'b101;
		y[592] = 12'b111111100010;
		z[592] = 3'b011;
		y[593] = 12'b001111111110;
		z[593] = 3'b110;
		y[594] = 12'b001111111111;
		z[594] = 3'b110;
		y[595] = 12'b010111101010;
		z[595] = 3'b111;
		y[596] = 12'b101110001010;
		z[596] = 3'b101;
		y[597] = 12'b101011001111;
		z[597] = 3'b101;
		y[598] = 12'b100101111011;
		z[598] = 3'b110;
		y[599] = 12'b000110000110;
		z[599] = 3'b000;
		y[600] = 12'b100001010100;
		z[600] = 3'b100;
		y[601] = 12'b110000011001;
		z[601] = 3'b001;
		y[602] = 12'b110110001010;
		z[602] = 3'b101;
		y[603] = 12'b010101001011;
		z[603] = 3'b010;
		y[604] = 12'b101011110100;
		z[604] = 3'b001;
		y[605] = 12'b000101111101;
		z[605] = 3'b111;
		y[606] = 12'b001101011101;
		z[606] = 3'b001;
		y[607] = 12'b111011101001;
		z[607] = 3'b110;
		y[608] = 12'b000111010110;
		z[608] = 3'b101;
		y[609] = 12'b101001000011;
		z[609] = 3'b000;
		y[610] = 12'b000100111000;
		z[610] = 3'b101;
		y[611] = 12'b010100100011;
		z[611] = 3'b101;
		y[612] = 12'b101000001010;
		z[612] = 3'b111;
		y[613] = 12'b101110101001;
		z[613] = 3'b001;
		y[614] = 12'b101001011100;
		z[614] = 3'b001;
		y[615] = 12'b110100101011;
		z[615] = 3'b011;
		y[616] = 12'b010010001100;
		z[616] = 3'b000;
		y[617] = 12'b001100101111;
		z[617] = 3'b110;
		y[618] = 12'b001000101010;
		z[618] = 3'b101;
		y[619] = 12'b010100110011;
		z[619] = 3'b011;
		y[620] = 12'b011110111010;
		z[620] = 3'b101;
		y[621] = 12'b000101010111;
		z[621] = 3'b010;
		y[622] = 12'b001100011010;
		z[622] = 3'b000;
		y[623] = 12'b111011010111;
		z[623] = 3'b000;
		y[624] = 12'b100111101100;
		z[624] = 3'b101;
		y[625] = 12'b111011010011;
		z[625] = 3'b010;
		y[626] = 12'b010000101001;
		z[626] = 3'b010;
		y[627] = 12'b001000110011;
		z[627] = 3'b010;
		y[628] = 12'b111111010011;
		z[628] = 3'b110;
		y[629] = 12'b011110111111;
		z[629] = 3'b101;
		y[630] = 12'b011010110001;
		z[630] = 3'b001;
		y[631] = 12'b001110100011;
		z[631] = 3'b001;
		y[632] = 12'b001100100001;
		z[632] = 3'b011;
		y[633] = 12'b111010101011;
		z[633] = 3'b100;
		y[634] = 12'b100101001000;
		z[634] = 3'b000;
		y[635] = 12'b100000011110;
		z[635] = 3'b110;
		y[636] = 12'b010100100110;
		z[636] = 3'b111;
		y[637] = 12'b111110111000;
		z[637] = 3'b111;
		y[638] = 12'b100111101110;
		z[638] = 3'b111;
		y[639] = 12'b111101100011;
		z[639] = 3'b000;
		y[640] = 12'b000101000000;
		z[640] = 3'b111;
		y[641] = 12'b010101111100;
		z[641] = 3'b101;
		y[642] = 12'b100101100000;
		z[642] = 3'b011;
		y[643] = 12'b011100100010;
		z[643] = 3'b111;
		y[644] = 12'b010100011101;
		z[644] = 3'b100;
		y[645] = 12'b101001001010;
		z[645] = 3'b111;
		y[646] = 12'b101010010000;
		z[646] = 3'b110;
		y[647] = 12'b010001010100;
		z[647] = 3'b101;
		y[648] = 12'b110110011111;
		z[648] = 3'b100;
		y[649] = 12'b010101011011;
		z[649] = 3'b100;
		y[650] = 12'b001001001100;
		z[650] = 3'b110;
		y[651] = 12'b101010101010;
		z[651] = 3'b111;
		y[652] = 12'b001101101111;
		z[652] = 3'b010;
		y[653] = 12'b001011110000;
		z[653] = 3'b001;
		y[654] = 12'b110001111111;
		z[654] = 3'b100;
		y[655] = 12'b110001110111;
		z[655] = 3'b100;
		y[656] = 12'b001010011010;
		z[656] = 3'b110;
		y[657] = 12'b010000111111;
		z[657] = 3'b110;
		y[658] = 12'b011110110000;
		z[658] = 3'b111;
		y[659] = 12'b110011010110;
		z[659] = 3'b001;
		y[660] = 12'b100100101111;
		z[660] = 3'b110;
		y[661] = 12'b101111110111;
		z[661] = 3'b010;
		y[662] = 12'b101111100001;
		z[662] = 3'b001;
		y[663] = 12'b110010000010;
		z[663] = 3'b100;
		y[664] = 12'b001110111010;
		z[664] = 3'b011;
		y[665] = 12'b000010001001;
		z[665] = 3'b100;
		y[666] = 12'b000000001010;
		z[666] = 3'b000;
		y[667] = 12'b101110100000;
		z[667] = 3'b111;
		y[668] = 12'b011110011101;
		z[668] = 3'b010;
		y[669] = 12'b100011010011;
		z[669] = 3'b101;
		y[670] = 12'b111101111010;
		z[670] = 3'b010;
		y[671] = 12'b010110100100;
		z[671] = 3'b101;
		y[672] = 12'b000010001111;
		z[672] = 3'b000;
		y[673] = 12'b111001000111;
		z[673] = 3'b111;
		y[674] = 12'b001110101000;
		z[674] = 3'b000;
		y[675] = 12'b111010010001;
		z[675] = 3'b011;
		y[676] = 12'b110011001000;
		z[676] = 3'b111;
		y[677] = 12'b110111010001;
		z[677] = 3'b101;
		y[678] = 12'b100101101111;
		z[678] = 3'b101;
		y[679] = 12'b110000011101;
		z[679] = 3'b111;
		y[680] = 12'b111111011011;
		z[680] = 3'b001;
		y[681] = 12'b100111100101;
		z[681] = 3'b001;
		y[682] = 12'b101010110101;
		z[682] = 3'b101;
		y[683] = 12'b010001011000;
		z[683] = 3'b110;
		y[684] = 12'b111000100011;
		z[684] = 3'b110;
		y[685] = 12'b011011001111;
		z[685] = 3'b001;
		y[686] = 12'b111000011011;
		z[686] = 3'b001;
		y[687] = 12'b011110011101;
		z[687] = 3'b111;
		y[688] = 12'b110001010001;
		z[688] = 3'b100;
		y[689] = 12'b010101111101;
		z[689] = 3'b101;
		y[690] = 12'b011100110100;
		z[690] = 3'b100;
		y[691] = 12'b111001101011;
		z[691] = 3'b011;
		y[692] = 12'b100110110111;
		z[692] = 3'b101;
		y[693] = 12'b111111101000;
		z[693] = 3'b010;
		y[694] = 12'b101000011100;
		z[694] = 3'b010;
		y[695] = 12'b001001000010;
		z[695] = 3'b000;
		y[696] = 12'b011100111100;
		z[696] = 3'b111;
		y[697] = 12'b001000100010;
		z[697] = 3'b111;
		y[698] = 12'b111011111101;
		z[698] = 3'b011;
		y[699] = 12'b000001101000;
		z[699] = 3'b010;
		y[700] = 12'b000011000001;
		z[700] = 3'b010;
		y[701] = 12'b010000110001;
		z[701] = 3'b110;
		y[702] = 12'b101000111001;
		z[702] = 3'b000;
		y[703] = 12'b011100101001;
		z[703] = 3'b001;
		y[704] = 12'b101101111011;
		z[704] = 3'b001;
		y[705] = 12'b101110100010;
		z[705] = 3'b011;
		y[706] = 12'b101100000110;
		z[706] = 3'b111;
		y[707] = 12'b001100001101;
		z[707] = 3'b101;
		y[708] = 12'b000000001001;
		z[708] = 3'b010;
		y[709] = 12'b001101010111;
		z[709] = 3'b101;
		y[710] = 12'b000001100010;
		z[710] = 3'b010;
		y[711] = 12'b110100100111;
		z[711] = 3'b001;
		y[712] = 12'b000000111100;
		z[712] = 3'b110;
		y[713] = 12'b100111111001;
		z[713] = 3'b110;
		y[714] = 12'b110011000010;
		z[714] = 3'b100;
		y[715] = 12'b101010101110;
		z[715] = 3'b111;
		y[716] = 12'b110011100010;
		z[716] = 3'b000;
		y[717] = 12'b111100010110;
		z[717] = 3'b010;
		y[718] = 12'b011000010011;
		z[718] = 3'b101;
		y[719] = 12'b100100011001;
		z[719] = 3'b001;
		y[720] = 12'b000001001111;
		z[720] = 3'b101;
		y[721] = 12'b000001110101;
		z[721] = 3'b000;
		y[722] = 12'b011111001010;
		z[722] = 3'b111;
		y[723] = 12'b110110100101;
		z[723] = 3'b010;
		y[724] = 12'b010100010111;
		z[724] = 3'b011;
		y[725] = 12'b001100101010;
		z[725] = 3'b010;
		y[726] = 12'b000000000111;
		z[726] = 3'b000;
		y[727] = 12'b111010010001;
		z[727] = 3'b110;
		y[728] = 12'b111101101000;
		z[728] = 3'b001;
		y[729] = 12'b110000000101;
		z[729] = 3'b110;
		y[730] = 12'b101101101101;
		z[730] = 3'b101;
		y[731] = 12'b101111011100;
		z[731] = 3'b111;
		y[732] = 12'b110001010100;
		z[732] = 3'b000;
		y[733] = 12'b110101100001;
		z[733] = 3'b101;
		y[734] = 12'b101010111100;
		z[734] = 3'b010;
		y[735] = 12'b111000001010;
		z[735] = 3'b101;
		y[736] = 12'b000101100011;
		z[736] = 3'b101;
		y[737] = 12'b101100111110;
		z[737] = 3'b110;
		y[738] = 12'b001111101100;
		z[738] = 3'b110;
		y[739] = 12'b010001100010;
		z[739] = 3'b111;
		y[740] = 12'b000101101111;
		z[740] = 3'b011;
		y[741] = 12'b111110111010;
		z[741] = 3'b010;
		y[742] = 12'b000101000100;
		z[742] = 3'b010;
		y[743] = 12'b100000010111;
		z[743] = 3'b111;
		y[744] = 12'b000101110100;
		z[744] = 3'b100;
		y[745] = 12'b000001010101;
		z[745] = 3'b000;
		y[746] = 12'b111100011110;
		z[746] = 3'b101;
		y[747] = 12'b000001001011;
		z[747] = 3'b100;
		y[748] = 12'b100010001010;
		z[748] = 3'b010;
		y[749] = 12'b100011000101;
		z[749] = 3'b111;
		y[750] = 12'b101111010000;
		z[750] = 3'b001;
		y[751] = 12'b010011000111;
		z[751] = 3'b111;
		y[752] = 12'b111011011111;
		z[752] = 3'b111;
		y[753] = 12'b011000011000;
		z[753] = 3'b101;
		y[754] = 12'b000000101110;
		z[754] = 3'b001;
		y[755] = 12'b100111111001;
		z[755] = 3'b110;
		y[756] = 12'b101101001011;
		z[756] = 3'b111;
		y[757] = 12'b100010101010;
		z[757] = 3'b111;
		y[758] = 12'b000010000110;
		z[758] = 3'b101;
		y[759] = 12'b010101001111;
		z[759] = 3'b010;
		y[760] = 12'b100010100001;
		z[760] = 3'b001;
		y[761] = 12'b001111100010;
		z[761] = 3'b010;
		y[762] = 12'b110010011011;
		z[762] = 3'b011;
		y[763] = 12'b000010010001;
		z[763] = 3'b100;
		y[764] = 12'b100010100000;
		z[764] = 3'b111;
		y[765] = 12'b101011111000;
		z[765] = 3'b010;
		y[766] = 12'b000001010110;
		z[766] = 3'b100;
		y[767] = 12'b010010101101;
		z[767] = 3'b011;
		y[768] = 12'b110111010010;
		z[768] = 3'b101;
		y[769] = 12'b011111000100;
		z[769] = 3'b101;
		y[770] = 12'b101110010111;
		z[770] = 3'b101;
		y[771] = 12'b010010010000;
		z[771] = 3'b101;
		y[772] = 12'b100001110000;
		z[772] = 3'b010;
		y[773] = 12'b110100100010;
		z[773] = 3'b100;
		y[774] = 12'b010001000010;
		z[774] = 3'b111;
		y[775] = 12'b101000011101;
		z[775] = 3'b011;
		y[776] = 12'b110010000001;
		z[776] = 3'b010;
		y[777] = 12'b101101110110;
		z[777] = 3'b001;
		y[778] = 12'b111101101001;
		z[778] = 3'b111;
		y[779] = 12'b000101001000;
		z[779] = 3'b111;
		y[780] = 12'b000101001011;
		z[780] = 3'b110;
		y[781] = 12'b011011011100;
		z[781] = 3'b001;
		y[782] = 12'b101011010000;
		z[782] = 3'b111;
		y[783] = 12'b001101110001;
		z[783] = 3'b101;
		y[784] = 12'b000011110101;
		z[784] = 3'b111;
		y[785] = 12'b111011011101;
		z[785] = 3'b101;
		y[786] = 12'b110000110110;
		z[786] = 3'b010;
		y[787] = 12'b110011011110;
		z[787] = 3'b110;
		y[788] = 12'b100001010101;
		z[788] = 3'b011;
		y[789] = 12'b001011000101;
		z[789] = 3'b101;
		y[790] = 12'b101100000011;
		z[790] = 3'b111;
		y[791] = 12'b101100000010;
		z[791] = 3'b000;
		y[792] = 12'b110010011100;
		z[792] = 3'b100;
		y[793] = 12'b111011011111;
		z[793] = 3'b100;
		y[794] = 12'b001111000100;
		z[794] = 3'b001;
		y[795] = 12'b000001000011;
		z[795] = 3'b110;
		y[796] = 12'b000010010101;
		z[796] = 3'b001;
		y[797] = 12'b011010011000;
		z[797] = 3'b100;
		y[798] = 12'b001100001001;
		z[798] = 3'b010;
		y[799] = 12'b111010011010;
		z[799] = 3'b010;
		y[800] = 12'b011111000011;
		z[800] = 3'b001;
		y[801] = 12'b001101001001;
		z[801] = 3'b100;
		y[802] = 12'b011110011100;
		z[802] = 3'b101;
		y[803] = 12'b100110000100;
		z[803] = 3'b110;
		y[804] = 12'b110010111001;
		z[804] = 3'b000;
		y[805] = 12'b110010000001;
		z[805] = 3'b000;
		y[806] = 12'b010001101001;
		z[806] = 3'b000;
		y[807] = 12'b110101110000;
		z[807] = 3'b100;
		y[808] = 12'b100011100001;
		z[808] = 3'b101;
		y[809] = 12'b000001101000;
		z[809] = 3'b101;
		y[810] = 12'b011010011110;
		z[810] = 3'b101;
		y[811] = 12'b011010100101;
		z[811] = 3'b000;
		y[812] = 12'b111000011011;
		z[812] = 3'b011;
		y[813] = 12'b110101000010;
		z[813] = 3'b101;
		y[814] = 12'b110011110001;
		z[814] = 3'b100;
		y[815] = 12'b111100100000;
		z[815] = 3'b111;
		y[816] = 12'b000011111101;
		z[816] = 3'b101;
		y[817] = 12'b111101111011;
		z[817] = 3'b111;
		y[818] = 12'b000110010101;
		z[818] = 3'b111;
		y[819] = 12'b010010000111;
		z[819] = 3'b010;
		y[820] = 12'b101111010110;
		z[820] = 3'b001;
		y[821] = 12'b110011101101;
		z[821] = 3'b101;
		y[822] = 12'b011111110100;
		z[822] = 3'b101;
		y[823] = 12'b000011100001;
		z[823] = 3'b111;
		y[824] = 12'b110001010011;
		z[824] = 3'b100;
		y[825] = 12'b001001101111;
		z[825] = 3'b001;
		y[826] = 12'b001010001001;
		z[826] = 3'b100;
		y[827] = 12'b101101000011;
		z[827] = 3'b011;
		y[828] = 12'b110100101000;
		z[828] = 3'b000;
		y[829] = 12'b000110101100;
		z[829] = 3'b111;
		y[830] = 12'b011000000100;
		z[830] = 3'b001;
		y[831] = 12'b010111100100;
		z[831] = 3'b000;
		y[832] = 12'b000010100110;
		z[832] = 3'b101;
		y[833] = 12'b011101011010;
		z[833] = 3'b001;
		y[834] = 12'b010100001011;
		z[834] = 3'b001;
		y[835] = 12'b101100010110;
		z[835] = 3'b110;
		y[836] = 12'b110101110000;
		z[836] = 3'b000;
		y[837] = 12'b101011010001;
		z[837] = 3'b001;
		y[838] = 12'b110110111100;
		z[838] = 3'b010;
		y[839] = 12'b111000110011;
		z[839] = 3'b100;
		y[840] = 12'b000010011100;
		z[840] = 3'b010;
		y[841] = 12'b010011100110;
		z[841] = 3'b111;
		y[842] = 12'b000110001101;
		z[842] = 3'b111;
		y[843] = 12'b111110101011;
		z[843] = 3'b011;
		y[844] = 12'b100100001111;
		z[844] = 3'b001;
		y[845] = 12'b101000100001;
		z[845] = 3'b101;
		y[846] = 12'b111110101110;
		z[846] = 3'b110;
		y[847] = 12'b101111111100;
		z[847] = 3'b110;
		y[848] = 12'b010110110000;
		z[848] = 3'b010;
		y[849] = 12'b100100011100;
		z[849] = 3'b111;
		y[850] = 12'b000001111110;
		z[850] = 3'b110;
		y[851] = 12'b111111011001;
		z[851] = 3'b001;
		y[852] = 12'b011100111001;
		z[852] = 3'b000;
		y[853] = 12'b111110010100;
		z[853] = 3'b110;
		y[854] = 12'b001000000000;
		z[854] = 3'b011;
		y[855] = 12'b001010110011;
		z[855] = 3'b010;
		y[856] = 12'b110110000001;
		z[856] = 3'b001;
		y[857] = 12'b000011100011;
		z[857] = 3'b011;
		y[858] = 12'b111001000110;
		z[858] = 3'b011;
		y[859] = 12'b101101101010;
		z[859] = 3'b000;
		y[860] = 12'b100111011000;
		z[860] = 3'b010;
		y[861] = 12'b000011100101;
		z[861] = 3'b010;
		y[862] = 12'b001011101101;
		z[862] = 3'b011;
		y[863] = 12'b000110011100;
		z[863] = 3'b100;
		y[864] = 12'b100001011000;
		z[864] = 3'b100;
		y[865] = 12'b010111111010;
		z[865] = 3'b111;
		y[866] = 12'b110101011111;
		z[866] = 3'b000;
		y[867] = 12'b100100010100;
		z[867] = 3'b001;
		y[868] = 12'b010011110100;
		z[868] = 3'b010;
		y[869] = 12'b110010100010;
		z[869] = 3'b101;
		y[870] = 12'b101000011101;
		z[870] = 3'b110;
		y[871] = 12'b010000000111;
		z[871] = 3'b101;
		y[872] = 12'b100011110111;
		z[872] = 3'b001;
		y[873] = 12'b001110111101;
		z[873] = 3'b010;
		y[874] = 12'b010111011011;
		z[874] = 3'b110;
		y[875] = 12'b011111011100;
		z[875] = 3'b010;
		y[876] = 12'b110000001001;
		z[876] = 3'b110;
		y[877] = 12'b110110011000;
		z[877] = 3'b010;
		y[878] = 12'b110111000111;
		z[878] = 3'b000;
		y[879] = 12'b000100001111;
		z[879] = 3'b101;
		y[880] = 12'b111111001111;
		z[880] = 3'b001;
		y[881] = 12'b011010110100;
		z[881] = 3'b101;
		y[882] = 12'b110011001101;
		z[882] = 3'b000;
		y[883] = 12'b110011011000;
		z[883] = 3'b100;
		y[884] = 12'b101101111100;
		z[884] = 3'b010;
		y[885] = 12'b010011011100;
		z[885] = 3'b111;
		y[886] = 12'b000010010010;
		z[886] = 3'b000;
		y[887] = 12'b110111101100;
		z[887] = 3'b110;
		y[888] = 12'b100100101010;
		z[888] = 3'b000;
		y[889] = 12'b100001101100;
		z[889] = 3'b111;
		y[890] = 12'b001001110011;
		z[890] = 3'b100;
		y[891] = 12'b101001100010;
		z[891] = 3'b011;
		y[892] = 12'b100101100011;
		z[892] = 3'b001;
		y[893] = 12'b111100001011;
		z[893] = 3'b101;
		y[894] = 12'b100010111010;
		z[894] = 3'b111;
		y[895] = 12'b000000011100;
		z[895] = 3'b000;
		y[896] = 12'b001100010110;
		z[896] = 3'b000;
		y[897] = 12'b111011010111;
		z[897] = 3'b110;
		y[898] = 12'b000010101010;
		z[898] = 3'b100;
		y[899] = 12'b110011001000;
		z[899] = 3'b001;
		y[900] = 12'b101000111111;
		z[900] = 3'b101;
		y[901] = 12'b111000001000;
		z[901] = 3'b110;
		y[902] = 12'b010101000110;
		z[902] = 3'b000;
		y[903] = 12'b101000110010;
		z[903] = 3'b101;
		y[904] = 12'b111001110011;
		z[904] = 3'b100;
		y[905] = 12'b111011101010;
		z[905] = 3'b100;
		y[906] = 12'b000000111111;
		z[906] = 3'b110;
		y[907] = 12'b100111010101;
		z[907] = 3'b111;
		y[908] = 12'b000010000000;
		z[908] = 3'b110;
		y[909] = 12'b110011010101;
		z[909] = 3'b100;
		y[910] = 12'b000010001110;
		z[910] = 3'b110;
		y[911] = 12'b011111000110;
		z[911] = 3'b010;
		y[912] = 12'b011001010111;
		z[912] = 3'b110;
		y[913] = 12'b011000001110;
		z[913] = 3'b001;
		y[914] = 12'b010111011001;
		z[914] = 3'b011;
		y[915] = 12'b001001000010;
		z[915] = 3'b100;
		y[916] = 12'b001000100101;
		z[916] = 3'b100;
		y[917] = 12'b001101010001;
		z[917] = 3'b000;
		y[918] = 12'b111111100100;
		z[918] = 3'b010;
		y[919] = 12'b011010000010;
		z[919] = 3'b110;
		y[920] = 12'b100000111101;
		z[920] = 3'b111;
		y[921] = 12'b101111011101;
		z[921] = 3'b100;
		y[922] = 12'b111001100111;
		z[922] = 3'b001;
		y[923] = 12'b110011100010;
		z[923] = 3'b011;
		y[924] = 12'b011011010010;
		z[924] = 3'b111;
		y[925] = 12'b110000000001;
		z[925] = 3'b110;
		y[926] = 12'b100011000100;
		z[926] = 3'b110;
		y[927] = 12'b000010110101;
		z[927] = 3'b101;
		y[928] = 12'b110000001011;
		z[928] = 3'b010;
		y[929] = 12'b101100000000;
		z[929] = 3'b110;
		y[930] = 12'b001010001100;
		z[930] = 3'b101;
		y[931] = 12'b001010110011;
		z[931] = 3'b101;
		y[932] = 12'b000000000101;
		z[932] = 3'b000;
		y[933] = 12'b010100101111;
		z[933] = 3'b011;
		y[934] = 12'b010100111001;
		z[934] = 3'b101;
		y[935] = 12'b100100111101;
		z[935] = 3'b101;
		y[936] = 12'b101101111001;
		z[936] = 3'b010;
		y[937] = 12'b101001001000;
		z[937] = 3'b010;
		y[938] = 12'b110110011111;
		z[938] = 3'b101;
		y[939] = 12'b100110011001;
		z[939] = 3'b101;
		y[940] = 12'b110000110110;
		z[940] = 3'b010;
		y[941] = 12'b010111000111;
		z[941] = 3'b010;
		y[942] = 12'b010001000100;
		z[942] = 3'b111;
		y[943] = 12'b111101101001;
		z[943] = 3'b100;
		y[944] = 12'b110101100010;
		z[944] = 3'b111;
		y[945] = 12'b111110011101;
		z[945] = 3'b010;
		y[946] = 12'b010011100110;
		z[946] = 3'b100;
		y[947] = 12'b001010011000;
		z[947] = 3'b010;
		y[948] = 12'b100101001110;
		z[948] = 3'b111;
		y[949] = 12'b111110110111;
		z[949] = 3'b001;
		y[950] = 12'b111010111101;
		z[950] = 3'b001;
		y[951] = 12'b111010010110;
		z[951] = 3'b010;
		y[952] = 12'b001001010101;
		z[952] = 3'b111;
		y[953] = 12'b010100001100;
		z[953] = 3'b101;
		y[954] = 12'b010000111010;
		z[954] = 3'b100;
		y[955] = 12'b100111101000;
		z[955] = 3'b111;
		y[956] = 12'b110101010111;
		z[956] = 3'b111;
		y[957] = 12'b100010011110;
		z[957] = 3'b010;
		y[958] = 12'b010000111110;
		z[958] = 3'b010;
		y[959] = 12'b100110111110;
		z[959] = 3'b101;
		y[960] = 12'b101110101001;
		z[960] = 3'b000;
		y[961] = 12'b101100010111;
		z[961] = 3'b101;
		y[962] = 12'b000110110110;
		z[962] = 3'b000;
		y[963] = 12'b010001001001;
		z[963] = 3'b010;
		y[964] = 12'b010000101110;
		z[964] = 3'b001;
		y[965] = 12'b011101001101;
		z[965] = 3'b001;
		y[966] = 12'b111001101011;
		z[966] = 3'b001;
		y[967] = 12'b010001011001;
		z[967] = 3'b110;
		y[968] = 12'b101100011101;
		z[968] = 3'b100;
		y[969] = 12'b110110111100;
		z[969] = 3'b101;
		y[970] = 12'b010100110010;
		z[970] = 3'b010;
		y[971] = 12'b101110110111;
		z[971] = 3'b001;
		y[972] = 12'b110001010111;
		z[972] = 3'b000;
		y[973] = 12'b101010111000;
		z[973] = 3'b111;
		y[974] = 12'b011111100111;
		z[974] = 3'b011;
		y[975] = 12'b110110001011;
		z[975] = 3'b111;
		y[976] = 12'b110001000101;
		z[976] = 3'b010;
		y[977] = 12'b000010111111;
		z[977] = 3'b100;
		y[978] = 12'b110010011010;
		z[978] = 3'b000;
		y[979] = 12'b011010000110;
		z[979] = 3'b101;
		y[980] = 12'b011001010111;
		z[980] = 3'b010;
		y[981] = 12'b110001000100;
		z[981] = 3'b110;
		y[982] = 12'b111111010101;
		z[982] = 3'b110;
		y[983] = 12'b010110100000;
		z[983] = 3'b111;
		y[984] = 12'b110011000000;
		z[984] = 3'b010;
		y[985] = 12'b101100100101;
		z[985] = 3'b001;
		y[986] = 12'b110001010010;
		z[986] = 3'b000;
		y[987] = 12'b001101001001;
		z[987] = 3'b011;
		y[988] = 12'b100010000110;
		z[988] = 3'b101;
		y[989] = 12'b100001000011;
		z[989] = 3'b000;
		y[990] = 12'b111110001111;
		z[990] = 3'b000;
		y[991] = 12'b111011001000;
		z[991] = 3'b110;
		y[992] = 12'b110110110100;
		z[992] = 3'b110;
		y[993] = 12'b101111110010;
		z[993] = 3'b101;
		y[994] = 12'b010110100101;
		z[994] = 3'b011;
		y[995] = 12'b101011101001;
		z[995] = 3'b101;
		y[996] = 12'b000001110011;
		z[996] = 3'b010;
		y[997] = 12'b100101111100;
		z[997] = 3'b100;
		y[998] = 12'b101001110111;
		z[998] = 3'b100;
		y[999] = 12'b010000011011;
		z[999] = 3'b110;
		y[1000] = 12'b000110110111;
		z[1000] = 3'b100;
		y[1001] = 12'b100110100100;
		z[1001] = 3'b100;
		y[1002] = 12'b001111111010;
		z[1002] = 3'b101;
		y[1003] = 12'b111010100010;
		z[1003] = 3'b011;
		y[1004] = 12'b100110011110;
		z[1004] = 3'b110;
		y[1005] = 12'b111010001111;
		z[1005] = 3'b001;
		y[1006] = 12'b100010101101;
		z[1006] = 3'b101;
		y[1007] = 12'b000010011000;
		z[1007] = 3'b101;
		y[1008] = 12'b101010110111;
		z[1008] = 3'b110;
		y[1009] = 12'b111111101010;
		z[1009] = 3'b111;
		y[1010] = 12'b111000101110;
		z[1010] = 3'b110;
		y[1011] = 12'b000000100011;
		z[1011] = 3'b001;
		y[1012] = 12'b101001001011;
		z[1012] = 3'b011;
		y[1013] = 12'b111100110110;
		z[1013] = 3'b000;
		y[1014] = 12'b111100000010;
		z[1014] = 3'b100;
		y[1015] = 12'b101001000011;
		z[1015] = 3'b110;
		y[1016] = 12'b011011110000;
		z[1016] = 3'b001;
		y[1017] = 12'b101100000111;
		z[1017] = 3'b101;
		y[1018] = 12'b110100000000;
		z[1018] = 3'b011;
		y[1019] = 12'b101101000100;
		z[1019] = 3'b101;
		y[1020] = 12'b001101001110;
		z[1020] = 3'b101;
		y[1021] = 12'b111101101011;
		z[1021] = 3'b001;
		y[1022] = 12'b101111111001;
		z[1022] = 3'b000;
		y[1023] = 12'b101111110111;
		z[1023] = 3'b101;
		y[1024] = 12'b001101001000;
		z[1024] = 3'b001;
		y[1025] = 12'b111101111001;
		z[1025] = 3'b000;
		y[1026] = 12'b110100001010;
		z[1026] = 3'b110;
		y[1027] = 12'b010000111000;
		z[1027] = 3'b010;
		y[1028] = 12'b000011101010;
		z[1028] = 3'b100;
		y[1029] = 12'b010100111000;
		z[1029] = 3'b101;
		y[1030] = 12'b111001110100;
		z[1030] = 3'b110;
		y[1031] = 12'b100111101101;
		z[1031] = 3'b011;
		y[1032] = 12'b101001001011;
		z[1032] = 3'b101;
		y[1033] = 12'b011100000100;
		z[1033] = 3'b011;
		y[1034] = 12'b011100001100;
		z[1034] = 3'b100;
		y[1035] = 12'b000010001101;
		z[1035] = 3'b110;
		y[1036] = 12'b111111111110;
		z[1036] = 3'b010;
		y[1037] = 12'b110000111000;
		z[1037] = 3'b011;
		y[1038] = 12'b001011101111;
		z[1038] = 3'b110;
		y[1039] = 12'b011010100011;
		z[1039] = 3'b010;
		y[1040] = 12'b111001011011;
		z[1040] = 3'b010;
		y[1041] = 12'b010111000111;
		z[1041] = 3'b010;
		y[1042] = 12'b110011111100;
		z[1042] = 3'b111;
		y[1043] = 12'b000011100011;
		z[1043] = 3'b111;
		y[1044] = 12'b011111011011;
		z[1044] = 3'b100;
		y[1045] = 12'b000111100011;
		z[1045] = 3'b110;
		y[1046] = 12'b110110110100;
		z[1046] = 3'b100;
		y[1047] = 12'b100011011011;
		z[1047] = 3'b100;
		y[1048] = 12'b011100100101;
		z[1048] = 3'b011;
		y[1049] = 12'b010011111001;
		z[1049] = 3'b010;
		y[1050] = 12'b111011000111;
		z[1050] = 3'b110;
		y[1051] = 12'b010001001111;
		z[1051] = 3'b000;
		y[1052] = 12'b100100010000;
		z[1052] = 3'b101;
		y[1053] = 12'b110101000010;
		z[1053] = 3'b011;
		y[1054] = 12'b000101100000;
		z[1054] = 3'b001;
		y[1055] = 12'b001010111111;
		z[1055] = 3'b000;
		y[1056] = 12'b001011001111;
		z[1056] = 3'b000;
		y[1057] = 12'b111000110000;
		z[1057] = 3'b010;
		y[1058] = 12'b110111000001;
		z[1058] = 3'b100;
		y[1059] = 12'b101101000101;
		z[1059] = 3'b111;
		y[1060] = 12'b000100000111;
		z[1060] = 3'b101;
		y[1061] = 12'b001000000000;
		z[1061] = 3'b000;
		y[1062] = 12'b111100110010;
		z[1062] = 3'b001;
		y[1063] = 12'b000110011011;
		z[1063] = 3'b111;
		y[1064] = 12'b101110110001;
		z[1064] = 3'b000;
		y[1065] = 12'b001101000001;
		z[1065] = 3'b011;
		y[1066] = 12'b110010010100;
		z[1066] = 3'b111;
		y[1067] = 12'b110100111000;
		z[1067] = 3'b110;
		y[1068] = 12'b101100110101;
		z[1068] = 3'b111;
		y[1069] = 12'b100010111000;
		z[1069] = 3'b111;
		y[1070] = 12'b001001101110;
		z[1070] = 3'b110;
		y[1071] = 12'b000110100100;
		z[1071] = 3'b101;
		y[1072] = 12'b101011011010;
		z[1072] = 3'b001;
		y[1073] = 12'b011001110101;
		z[1073] = 3'b010;
		y[1074] = 12'b110110000100;
		z[1074] = 3'b010;
		y[1075] = 12'b011100010101;
		z[1075] = 3'b111;
		y[1076] = 12'b000111000111;
		z[1076] = 3'b011;
		y[1077] = 12'b101010001001;
		z[1077] = 3'b100;
		y[1078] = 12'b001100001010;
		z[1078] = 3'b111;
		y[1079] = 12'b111111100000;
		z[1079] = 3'b110;
		y[1080] = 12'b010101110011;
		z[1080] = 3'b001;
		y[1081] = 12'b011001011111;
		z[1081] = 3'b100;
		y[1082] = 12'b100011000111;
		z[1082] = 3'b100;
		y[1083] = 12'b011000010111;
		z[1083] = 3'b001;
		y[1084] = 12'b100001001111;
		z[1084] = 3'b111;
		y[1085] = 12'b110000110000;
		z[1085] = 3'b110;
		y[1086] = 12'b101011100010;
		z[1086] = 3'b010;
		y[1087] = 12'b101101100101;
		z[1087] = 3'b001;
		y[1088] = 12'b100010110001;
		z[1088] = 3'b110;
		y[1089] = 12'b100000011100;
		z[1089] = 3'b100;
		y[1090] = 12'b000001111000;
		z[1090] = 3'b110;
		y[1091] = 12'b100000101101;
		z[1091] = 3'b000;
		y[1092] = 12'b100101010111;
		z[1092] = 3'b010;
		y[1093] = 12'b000001001100;
		z[1093] = 3'b011;
		y[1094] = 12'b001111100100;
		z[1094] = 3'b101;
		y[1095] = 12'b010100000100;
		z[1095] = 3'b000;
		y[1096] = 12'b000100001011;
		z[1096] = 3'b011;
		y[1097] = 12'b000110000010;
		z[1097] = 3'b001;
		y[1098] = 12'b000111110101;
		z[1098] = 3'b010;
		y[1099] = 12'b010101100000;
		z[1099] = 3'b011;
		y[1100] = 12'b000010111001;
		z[1100] = 3'b000;
		y[1101] = 12'b011110001101;
		z[1101] = 3'b010;
		y[1102] = 12'b010000011001;
		z[1102] = 3'b110;
		y[1103] = 12'b001011110010;
		z[1103] = 3'b000;
		y[1104] = 12'b010111000100;
		z[1104] = 3'b111;
		y[1105] = 12'b111100100011;
		z[1105] = 3'b101;
		y[1106] = 12'b010101010011;
		z[1106] = 3'b111;
		y[1107] = 12'b101010110011;
		z[1107] = 3'b110;
		y[1108] = 12'b110000110110;
		z[1108] = 3'b000;
		y[1109] = 12'b010111001000;
		z[1109] = 3'b001;
		y[1110] = 12'b101101001100;
		z[1110] = 3'b100;
		y[1111] = 12'b001111000011;
		z[1111] = 3'b001;
		y[1112] = 12'b010001110111;
		z[1112] = 3'b001;
		y[1113] = 12'b000001110100;
		z[1113] = 3'b000;
		y[1114] = 12'b101011110101;
		z[1114] = 3'b010;
		y[1115] = 12'b101000100101;
		z[1115] = 3'b100;
		y[1116] = 12'b011101110001;
		z[1116] = 3'b000;
		y[1117] = 12'b111001011101;
		z[1117] = 3'b001;
		y[1118] = 12'b010001000110;
		z[1118] = 3'b010;
		y[1119] = 12'b110111000000;
		z[1119] = 3'b110;
		y[1120] = 12'b110010110001;
		z[1120] = 3'b000;
		y[1121] = 12'b001011011010;
		z[1121] = 3'b011;
		y[1122] = 12'b001011010010;
		z[1122] = 3'b111;
		y[1123] = 12'b100101100010;
		z[1123] = 3'b110;
		y[1124] = 12'b011111011000;
		z[1124] = 3'b011;
		y[1125] = 12'b101010001100;
		z[1125] = 3'b000;
		y[1126] = 12'b010110011010;
		z[1126] = 3'b000;
		y[1127] = 12'b100100010011;
		z[1127] = 3'b010;
		y[1128] = 12'b010001001100;
		z[1128] = 3'b000;
		y[1129] = 12'b000010110010;
		z[1129] = 3'b001;
		y[1130] = 12'b111111111000;
		z[1130] = 3'b001;
		y[1131] = 12'b010010010001;
		z[1131] = 3'b011;
		y[1132] = 12'b100000000110;
		z[1132] = 3'b001;
		y[1133] = 12'b001111101101;
		z[1133] = 3'b001;
		y[1134] = 12'b010110110101;
		z[1134] = 3'b110;
		y[1135] = 12'b111100010001;
		z[1135] = 3'b110;
		y[1136] = 12'b110001000011;
		z[1136] = 3'b011;
		y[1137] = 12'b101001001100;
		z[1137] = 3'b100;
		y[1138] = 12'b100101110010;
		z[1138] = 3'b001;
		y[1139] = 12'b010110100110;
		z[1139] = 3'b011;
		y[1140] = 12'b110110010111;
		z[1140] = 3'b011;
		y[1141] = 12'b100001101011;
		z[1141] = 3'b001;
		y[1142] = 12'b000001001111;
		z[1142] = 3'b110;
		y[1143] = 12'b000100100000;
		z[1143] = 3'b011;
		y[1144] = 12'b011001101000;
		z[1144] = 3'b010;
		y[1145] = 12'b011101011010;
		z[1145] = 3'b111;
		y[1146] = 12'b001010000101;
		z[1146] = 3'b011;
		y[1147] = 12'b000011000110;
		z[1147] = 3'b010;
		y[1148] = 12'b001101011010;
		z[1148] = 3'b101;
		y[1149] = 12'b010110111011;
		z[1149] = 3'b001;
		y[1150] = 12'b001111101111;
		z[1150] = 3'b100;
		y[1151] = 12'b001101101000;
		z[1151] = 3'b111;
		y[1152] = 12'b101010000010;
		z[1152] = 3'b101;
		y[1153] = 12'b101001011110;
		z[1153] = 3'b001;
		y[1154] = 12'b101000111101;
		z[1154] = 3'b100;
		y[1155] = 12'b100000100100;
		z[1155] = 3'b111;
		y[1156] = 12'b100001010011;
		z[1156] = 3'b111;
		y[1157] = 12'b000000000010;
		z[1157] = 3'b111;
		y[1158] = 12'b000000110110;
		z[1158] = 3'b101;
		y[1159] = 12'b000001101110;
		z[1159] = 3'b100;
		y[1160] = 12'b101010001110;
		z[1160] = 3'b101;
		y[1161] = 12'b111010011110;
		z[1161] = 3'b100;
		y[1162] = 12'b111001000100;
		z[1162] = 3'b111;
		y[1163] = 12'b000101001100;
		z[1163] = 3'b100;
		y[1164] = 12'b001001011010;
		z[1164] = 3'b101;
		y[1165] = 12'b011001101010;
		z[1165] = 3'b010;
		y[1166] = 12'b000100101111;
		z[1166] = 3'b010;
		y[1167] = 12'b110110001111;
		z[1167] = 3'b110;
		y[1168] = 12'b111001111101;
		z[1168] = 3'b001;
		y[1169] = 12'b010011011101;
		z[1169] = 3'b110;
		y[1170] = 12'b011011100010;
		z[1170] = 3'b000;
		y[1171] = 12'b011101011101;
		z[1171] = 3'b011;
		y[1172] = 12'b101011000011;
		z[1172] = 3'b000;
		y[1173] = 12'b100101011101;
		z[1173] = 3'b000;
		y[1174] = 12'b111000101101;
		z[1174] = 3'b011;
		y[1175] = 12'b010100111110;
		z[1175] = 3'b000;
		y[1176] = 12'b011101001111;
		z[1176] = 3'b011;
		y[1177] = 12'b100000110101;
		z[1177] = 3'b101;
		y[1178] = 12'b101110111111;
		z[1178] = 3'b101;
		y[1179] = 12'b101000001010;
		z[1179] = 3'b111;
		y[1180] = 12'b011111100001;
		z[1180] = 3'b010;
		y[1181] = 12'b100110110100;
		z[1181] = 3'b011;
		y[1182] = 12'b000000011000;
		z[1182] = 3'b110;
		y[1183] = 12'b011110011100;
		z[1183] = 3'b100;
		y[1184] = 12'b000100011000;
		z[1184] = 3'b000;
		y[1185] = 12'b111000001111;
		z[1185] = 3'b010;
		y[1186] = 12'b001111100000;
		z[1186] = 3'b101;
		y[1187] = 12'b110011101110;
		z[1187] = 3'b000;
		y[1188] = 12'b100101011010;
		z[1188] = 3'b111;
		y[1189] = 12'b000101110111;
		z[1189] = 3'b100;
		y[1190] = 12'b011000101001;
		z[1190] = 3'b000;
		y[1191] = 12'b101100001011;
		z[1191] = 3'b011;
		y[1192] = 12'b011000011000;
		z[1192] = 3'b011;
		y[1193] = 12'b010001000010;
		z[1193] = 3'b001;
		y[1194] = 12'b101001010000;
		z[1194] = 3'b110;
		y[1195] = 12'b010100001001;
		z[1195] = 3'b001;
		y[1196] = 12'b110101011011;
		z[1196] = 3'b010;
		y[1197] = 12'b101010111101;
		z[1197] = 3'b101;
		y[1198] = 12'b101010101111;
		z[1198] = 3'b000;
		y[1199] = 12'b000100001110;
		z[1199] = 3'b001;
		y[1200] = 12'b101001000100;
		z[1200] = 3'b110;
		y[1201] = 12'b010011001101;
		z[1201] = 3'b000;
		y[1202] = 12'b010110110011;
		z[1202] = 3'b110;
		y[1203] = 12'b011000001001;
		z[1203] = 3'b101;
		y[1204] = 12'b010101010011;
		z[1204] = 3'b101;
		y[1205] = 12'b000011001000;
		z[1205] = 3'b100;
		y[1206] = 12'b100001000000;
		z[1206] = 3'b100;
		y[1207] = 12'b100000101010;
		z[1207] = 3'b001;
		y[1208] = 12'b001110101001;
		z[1208] = 3'b000;
		y[1209] = 12'b000100000001;
		z[1209] = 3'b101;
		y[1210] = 12'b111011111110;
		z[1210] = 3'b101;
		y[1211] = 12'b010101111100;
		z[1211] = 3'b000;
		y[1212] = 12'b010001110001;
		z[1212] = 3'b100;
		y[1213] = 12'b011101011100;
		z[1213] = 3'b100;
		y[1214] = 12'b011101010111;
		z[1214] = 3'b110;
		y[1215] = 12'b100111010100;
		z[1215] = 3'b001;
		y[1216] = 12'b010011111101;
		z[1216] = 3'b000;
		y[1217] = 12'b010101100111;
		z[1217] = 3'b000;
		y[1218] = 12'b110001000110;
		z[1218] = 3'b010;
		y[1219] = 12'b111001010000;
		z[1219] = 3'b111;
		y[1220] = 12'b101001011111;
		z[1220] = 3'b010;
		y[1221] = 12'b000000100001;
		z[1221] = 3'b100;
		y[1222] = 12'b010001001010;
		z[1222] = 3'b011;
		y[1223] = 12'b000110111100;
		z[1223] = 3'b000;
		y[1224] = 12'b100001010010;
		z[1224] = 3'b110;
		y[1225] = 12'b000101111000;
		z[1225] = 3'b100;
		y[1226] = 12'b100101111110;
		z[1226] = 3'b101;
		y[1227] = 12'b100010010011;
		z[1227] = 3'b100;
		y[1228] = 12'b110011000010;
		z[1228] = 3'b001;
		y[1229] = 12'b101111101110;
		z[1229] = 3'b000;
		y[1230] = 12'b111010001101;
		z[1230] = 3'b111;
		y[1231] = 12'b011011001111;
		z[1231] = 3'b101;
		y[1232] = 12'b000110111101;
		z[1232] = 3'b001;
		y[1233] = 12'b110101010011;
		z[1233] = 3'b110;
		y[1234] = 12'b011101011011;
		z[1234] = 3'b010;
		y[1235] = 12'b011110100110;
		z[1235] = 3'b110;
		y[1236] = 12'b010101000111;
		z[1236] = 3'b111;
		y[1237] = 12'b100110100110;
		z[1237] = 3'b101;
		y[1238] = 12'b101101101100;
		z[1238] = 3'b110;
		y[1239] = 12'b110101100010;
		z[1239] = 3'b001;
		y[1240] = 12'b000111000000;
		z[1240] = 3'b011;
		y[1241] = 12'b001111110110;
		z[1241] = 3'b010;
		y[1242] = 12'b111100110110;
		z[1242] = 3'b011;
		y[1243] = 12'b101101100001;
		z[1243] = 3'b111;
		y[1244] = 12'b011011000111;
		z[1244] = 3'b100;
		y[1245] = 12'b100110001100;
		z[1245] = 3'b101;
		y[1246] = 12'b111110011010;
		z[1246] = 3'b100;
		y[1247] = 12'b110111101011;
		z[1247] = 3'b010;
		y[1248] = 12'b111011100011;
		z[1248] = 3'b001;
		y[1249] = 12'b010110001010;
		z[1249] = 3'b100;
		y[1250] = 12'b100100111101;
		z[1250] = 3'b011;
		y[1251] = 12'b000001000110;
		z[1251] = 3'b011;
		y[1252] = 12'b100011000011;
		z[1252] = 3'b010;
		y[1253] = 12'b011110001110;
		z[1253] = 3'b101;
		y[1254] = 12'b111000001110;
		z[1254] = 3'b101;
		y[1255] = 12'b011001100110;
		z[1255] = 3'b100;
		y[1256] = 12'b001010101111;
		z[1256] = 3'b111;
		y[1257] = 12'b111111001100;
		z[1257] = 3'b000;
		y[1258] = 12'b000000111001;
		z[1258] = 3'b010;
		y[1259] = 12'b110101010010;
		z[1259] = 3'b100;
		y[1260] = 12'b010000101101;
		z[1260] = 3'b000;
		y[1261] = 12'b010000011101;
		z[1261] = 3'b010;
		y[1262] = 12'b101101110111;
		z[1262] = 3'b001;
		y[1263] = 12'b100110001000;
		z[1263] = 3'b000;
		y[1264] = 12'b001011111101;
		z[1264] = 3'b110;
		y[1265] = 12'b110110000011;
		z[1265] = 3'b011;
		y[1266] = 12'b001011011110;
		z[1266] = 3'b111;
		y[1267] = 12'b010010001100;
		z[1267] = 3'b110;
		y[1268] = 12'b001111101011;
		z[1268] = 3'b110;
		y[1269] = 12'b010000010101;
		z[1269] = 3'b100;
		y[1270] = 12'b011110010100;
		z[1270] = 3'b100;
		y[1271] = 12'b011000011111;
		z[1271] = 3'b101;
		y[1272] = 12'b111101101011;
		z[1272] = 3'b010;
		y[1273] = 12'b101110110010;
		z[1273] = 3'b000;
		y[1274] = 12'b011000101001;
		z[1274] = 3'b101;
		y[1275] = 12'b110011010100;
		z[1275] = 3'b100;
		y[1276] = 12'b111011011110;
		z[1276] = 3'b100;
		y[1277] = 12'b000000100110;
		z[1277] = 3'b001;
		y[1278] = 12'b000101010001;
		z[1278] = 3'b100;
		y[1279] = 12'b000111101011;
		z[1279] = 3'b101;
		y[1280] = 12'b000011011101;
		z[1280] = 3'b010;
		y[1281] = 12'b100100010010;
		z[1281] = 3'b001;
		y[1282] = 12'b110011110001;
		z[1282] = 3'b101;
		y[1283] = 12'b110100111101;
		z[1283] = 3'b000;
		y[1284] = 12'b101110010000;
		z[1284] = 3'b100;
		y[1285] = 12'b001000001101;
		z[1285] = 3'b101;
		y[1286] = 12'b101100101001;
		z[1286] = 3'b011;
		y[1287] = 12'b110111011110;
		z[1287] = 3'b010;
		y[1288] = 12'b100001011101;
		z[1288] = 3'b110;
		y[1289] = 12'b001010011100;
		z[1289] = 3'b010;
		y[1290] = 12'b100100000100;
		z[1290] = 3'b001;
		y[1291] = 12'b100010111000;
		z[1291] = 3'b010;
		y[1292] = 12'b001111101000;
		z[1292] = 3'b001;
		y[1293] = 12'b001000100011;
		z[1293] = 3'b000;
		y[1294] = 12'b110011010110;
		z[1294] = 3'b000;
		y[1295] = 12'b110100001111;
		z[1295] = 3'b000;
		y[1296] = 12'b110100110011;
		z[1296] = 3'b100;
		y[1297] = 12'b101011100001;
		z[1297] = 3'b010;
		y[1298] = 12'b100101101110;
		z[1298] = 3'b010;
		y[1299] = 12'b111101110010;
		z[1299] = 3'b011;
		y[1300] = 12'b011011111100;
		z[1300] = 3'b110;
		y[1301] = 12'b011000110100;
		z[1301] = 3'b101;
		y[1302] = 12'b001001000100;
		z[1302] = 3'b010;
		y[1303] = 12'b101101111011;
		z[1303] = 3'b011;
		y[1304] = 12'b100010110101;
		z[1304] = 3'b011;
		y[1305] = 12'b011110011010;
		z[1305] = 3'b100;
		y[1306] = 12'b011000000011;
		z[1306] = 3'b000;
		y[1307] = 12'b101010011100;
		z[1307] = 3'b101;
		y[1308] = 12'b011010001110;
		z[1308] = 3'b110;
		y[1309] = 12'b111010100000;
		z[1309] = 3'b010;
		y[1310] = 12'b001000010111;
		z[1310] = 3'b110;
		y[1311] = 12'b011010100101;
		z[1311] = 3'b011;
		y[1312] = 12'b100001101011;
		z[1312] = 3'b001;
		y[1313] = 12'b111001100110;
		z[1313] = 3'b011;
		y[1314] = 12'b011110001000;
		z[1314] = 3'b111;
		y[1315] = 12'b110001011001;
		z[1315] = 3'b010;
		y[1316] = 12'b100111101010;
		z[1316] = 3'b010;
		y[1317] = 12'b011000111011;
		z[1317] = 3'b001;
		y[1318] = 12'b000010111001;
		z[1318] = 3'b001;
		y[1319] = 12'b000011100100;
		z[1319] = 3'b111;
		y[1320] = 12'b001011110011;
		z[1320] = 3'b001;
		y[1321] = 12'b111100001010;
		z[1321] = 3'b111;
		y[1322] = 12'b101001000101;
		z[1322] = 3'b011;
		y[1323] = 12'b101101011000;
		z[1323] = 3'b000;
		y[1324] = 12'b011011010001;
		z[1324] = 3'b110;
		y[1325] = 12'b001100100110;
		z[1325] = 3'b001;
		y[1326] = 12'b111111001111;
		z[1326] = 3'b100;
		y[1327] = 12'b111101111101;
		z[1327] = 3'b010;
		y[1328] = 12'b110111000011;
		z[1328] = 3'b001;
		y[1329] = 12'b100111000010;
		z[1329] = 3'b101;
		y[1330] = 12'b101011011101;
		z[1330] = 3'b001;
		y[1331] = 12'b010011000011;
		z[1331] = 3'b110;
		y[1332] = 12'b101101110111;
		z[1332] = 3'b001;
		y[1333] = 12'b011111001011;
		z[1333] = 3'b010;
		y[1334] = 12'b100111111011;
		z[1334] = 3'b010;
		y[1335] = 12'b110100100101;
		z[1335] = 3'b011;
		y[1336] = 12'b001000111001;
		z[1336] = 3'b000;
		y[1337] = 12'b110111000101;
		z[1337] = 3'b010;
		y[1338] = 12'b000010110010;
		z[1338] = 3'b101;
		y[1339] = 12'b010001000000;
		z[1339] = 3'b110;
		y[1340] = 12'b111011111001;
		z[1340] = 3'b001;
		y[1341] = 12'b100100111001;
		z[1341] = 3'b111;
		y[1342] = 12'b001111010101;
		z[1342] = 3'b011;
		y[1343] = 12'b001011000010;
		z[1343] = 3'b001;
		y[1344] = 12'b100000100111;
		z[1344] = 3'b111;
		y[1345] = 12'b010011110100;
		z[1345] = 3'b100;
		y[1346] = 12'b100100111111;
		z[1346] = 3'b100;
		y[1347] = 12'b011000010000;
		z[1347] = 3'b101;
		y[1348] = 12'b100011110101;
		z[1348] = 3'b011;
		y[1349] = 12'b010001110111;
		z[1349] = 3'b011;
		y[1350] = 12'b010100100101;
		z[1350] = 3'b001;
		y[1351] = 12'b000110110100;
		z[1351] = 3'b100;
		y[1352] = 12'b001010111100;
		z[1352] = 3'b001;
		y[1353] = 12'b011110100100;
		z[1353] = 3'b001;
		y[1354] = 12'b101101001100;
		z[1354] = 3'b001;
		y[1355] = 12'b000010101101;
		z[1355] = 3'b101;
		y[1356] = 12'b011111011001;
		z[1356] = 3'b000;
		y[1357] = 12'b111001100100;
		z[1357] = 3'b100;
		y[1358] = 12'b010110011110;
		z[1358] = 3'b111;
		y[1359] = 12'b000100110111;
		z[1359] = 3'b010;
		y[1360] = 12'b100101011100;
		z[1360] = 3'b101;
		y[1361] = 12'b111010100111;
		z[1361] = 3'b011;
		y[1362] = 12'b101100110101;
		z[1362] = 3'b011;
		y[1363] = 12'b010100001010;
		z[1363] = 3'b001;
		y[1364] = 12'b001001011001;
		z[1364] = 3'b100;
		y[1365] = 12'b000000011001;
		z[1365] = 3'b011;
		y[1366] = 12'b111100111101;
		z[1366] = 3'b001;
		y[1367] = 12'b100101010100;
		z[1367] = 3'b101;
		y[1368] = 12'b001010111011;
		z[1368] = 3'b000;
		y[1369] = 12'b111000110010;
		z[1369] = 3'b011;
		y[1370] = 12'b101101000000;
		z[1370] = 3'b001;
		y[1371] = 12'b110111011000;
		z[1371] = 3'b001;
		y[1372] = 12'b110111111111;
		z[1372] = 3'b000;
		y[1373] = 12'b111110110111;
		z[1373] = 3'b001;
		y[1374] = 12'b000001001011;
		z[1374] = 3'b010;
		y[1375] = 12'b110100011010;
		z[1375] = 3'b100;
		y[1376] = 12'b100001110111;
		z[1376] = 3'b100;
		y[1377] = 12'b100111110010;
		z[1377] = 3'b100;
		y[1378] = 12'b101110001101;
		z[1378] = 3'b110;
		y[1379] = 12'b100100101000;
		z[1379] = 3'b111;
		y[1380] = 12'b101100101111;
		z[1380] = 3'b101;
		y[1381] = 12'b001011100111;
		z[1381] = 3'b100;
		y[1382] = 12'b011111011001;
		z[1382] = 3'b010;
		y[1383] = 12'b110111010100;
		z[1383] = 3'b110;
		y[1384] = 12'b010011010001;
		z[1384] = 3'b111;
		y[1385] = 12'b010010011110;
		z[1385] = 3'b100;
		y[1386] = 12'b100010110011;
		z[1386] = 3'b010;
		y[1387] = 12'b110000000010;
		z[1387] = 3'b111;
		y[1388] = 12'b000001110110;
		z[1388] = 3'b111;
		y[1389] = 12'b101010010110;
		z[1389] = 3'b011;
		y[1390] = 12'b110001110001;
		z[1390] = 3'b001;
		y[1391] = 12'b100100100110;
		z[1391] = 3'b111;
		y[1392] = 12'b010111010100;
		z[1392] = 3'b011;
		y[1393] = 12'b011101001011;
		z[1393] = 3'b000;
		y[1394] = 12'b010110101111;
		z[1394] = 3'b111;
		y[1395] = 12'b101000110101;
		z[1395] = 3'b110;
		y[1396] = 12'b000000100111;
		z[1396] = 3'b011;
		y[1397] = 12'b001001101100;
		z[1397] = 3'b011;
		y[1398] = 12'b100000000101;
		z[1398] = 3'b101;
		y[1399] = 12'b010010110011;
		z[1399] = 3'b111;
		y[1400] = 12'b000111011001;
		z[1400] = 3'b011;
		y[1401] = 12'b011000110011;
		z[1401] = 3'b110;
		y[1402] = 12'b001001000111;
		z[1402] = 3'b100;
		y[1403] = 12'b011110001011;
		z[1403] = 3'b111;
		y[1404] = 12'b001110100000;
		z[1404] = 3'b010;
		y[1405] = 12'b101001001110;
		z[1405] = 3'b001;
		y[1406] = 12'b101010000110;
		z[1406] = 3'b001;
		y[1407] = 12'b111110000111;
		z[1407] = 3'b000;
		y[1408] = 12'b001101010110;
		z[1408] = 3'b100;
		y[1409] = 12'b100000100110;
		z[1409] = 3'b011;
		y[1410] = 12'b101110101101;
		z[1410] = 3'b000;
		y[1411] = 12'b010011011111;
		z[1411] = 3'b101;
		y[1412] = 12'b111101000000;
		z[1412] = 3'b011;
		y[1413] = 12'b000101010101;
		z[1413] = 3'b010;
		y[1414] = 12'b000011101010;
		z[1414] = 3'b111;
		y[1415] = 12'b010100111101;
		z[1415] = 3'b100;
		y[1416] = 12'b000000100100;
		z[1416] = 3'b110;
		y[1417] = 12'b011010011000;
		z[1417] = 3'b101;
		y[1418] = 12'b110110011000;
		z[1418] = 3'b111;
		y[1419] = 12'b110111010010;
		z[1419] = 3'b011;
		y[1420] = 12'b111110010010;
		z[1420] = 3'b100;
		y[1421] = 12'b001101111101;
		z[1421] = 3'b111;
		y[1422] = 12'b000110111011;
		z[1422] = 3'b111;
		y[1423] = 12'b010101100110;
		z[1423] = 3'b111;
		y[1424] = 12'b100111100110;
		z[1424] = 3'b100;
		y[1425] = 12'b011010001001;
		z[1425] = 3'b010;
		y[1426] = 12'b010011101001;
		z[1426] = 3'b110;
		y[1427] = 12'b100011110111;
		z[1427] = 3'b101;
		y[1428] = 12'b100110011110;
		z[1428] = 3'b010;
		y[1429] = 12'b110001101001;
		z[1429] = 3'b100;
		y[1430] = 12'b110010010111;
		z[1430] = 3'b101;
		y[1431] = 12'b100000010000;
		z[1431] = 3'b101;
		y[1432] = 12'b101101111010;
		z[1432] = 3'b011;
		y[1433] = 12'b001000111110;
		z[1433] = 3'b111;
		y[1434] = 12'b011011110001;
		z[1434] = 3'b001;
		y[1435] = 12'b011101001111;
		z[1435] = 3'b111;
		y[1436] = 12'b010011001011;
		z[1436] = 3'b111;
		y[1437] = 12'b110110100011;
		z[1437] = 3'b000;
		y[1438] = 12'b101000011101;
		z[1438] = 3'b100;
		y[1439] = 12'b101111100011;
		z[1439] = 3'b101;
		y[1440] = 12'b101101100001;
		z[1440] = 3'b000;
		y[1441] = 12'b000110000101;
		z[1441] = 3'b111;
		y[1442] = 12'b111100010101;
		z[1442] = 3'b110;
		y[1443] = 12'b100000100101;
		z[1443] = 3'b011;
		y[1444] = 12'b110111001110;
		z[1444] = 3'b100;
		y[1445] = 12'b000010101010;
		z[1445] = 3'b011;
		y[1446] = 12'b110111100000;
		z[1446] = 3'b110;
		y[1447] = 12'b111000111111;
		z[1447] = 3'b111;
		y[1448] = 12'b010001101111;
		z[1448] = 3'b101;
		y[1449] = 12'b001111000101;
		z[1449] = 3'b000;
		y[1450] = 12'b001101110100;
		z[1450] = 3'b111;
		y[1451] = 12'b111000011110;
		z[1451] = 3'b000;
		y[1452] = 12'b011100000010;
		z[1452] = 3'b101;
		y[1453] = 12'b100100111011;
		z[1453] = 3'b100;
		y[1454] = 12'b111010101001;
		z[1454] = 3'b111;
		y[1455] = 12'b100000111100;
		z[1455] = 3'b001;
		y[1456] = 12'b001000000110;
		z[1456] = 3'b101;
		y[1457] = 12'b001000111110;
		z[1457] = 3'b001;
		y[1458] = 12'b100011110111;
		z[1458] = 3'b101;
		y[1459] = 12'b000100011101;
		z[1459] = 3'b101;
		y[1460] = 12'b011011100111;
		z[1460] = 3'b010;
		y[1461] = 12'b101010001110;
		z[1461] = 3'b101;
		y[1462] = 12'b100110101111;
		z[1462] = 3'b100;
		y[1463] = 12'b100000110000;
		z[1463] = 3'b110;
		y[1464] = 12'b011100000001;
		z[1464] = 3'b100;
		y[1465] = 12'b000101100010;
		z[1465] = 3'b101;
		y[1466] = 12'b110011101000;
		z[1466] = 3'b000;
		y[1467] = 12'b101100111001;
		z[1467] = 3'b111;
		y[1468] = 12'b101010001101;
		z[1468] = 3'b100;
		y[1469] = 12'b110110010110;
		z[1469] = 3'b011;
		y[1470] = 12'b010111110011;
		z[1470] = 3'b110;
		y[1471] = 12'b000100101000;
		z[1471] = 3'b011;
		y[1472] = 12'b111011010111;
		z[1472] = 3'b100;
		y[1473] = 12'b001100010001;
		z[1473] = 3'b111;
		y[1474] = 12'b001001101001;
		z[1474] = 3'b001;
		y[1475] = 12'b110100001111;
		z[1475] = 3'b101;
		y[1476] = 12'b010100000011;
		z[1476] = 3'b001;
		y[1477] = 12'b010110100000;
		z[1477] = 3'b000;
		y[1478] = 12'b010011100001;
		z[1478] = 3'b111;
		y[1479] = 12'b010100111010;
		z[1479] = 3'b011;
		y[1480] = 12'b001110101101;
		z[1480] = 3'b110;
		y[1481] = 12'b100110110010;
		z[1481] = 3'b000;
		y[1482] = 12'b010100111010;
		z[1482] = 3'b111;
		y[1483] = 12'b101000100011;
		z[1483] = 3'b010;
		y[1484] = 12'b011010101010;
		z[1484] = 3'b111;
		y[1485] = 12'b001010011001;
		z[1485] = 3'b000;
		y[1486] = 12'b100010001101;
		z[1486] = 3'b111;
		y[1487] = 12'b011010110000;
		z[1487] = 3'b100;
		y[1488] = 12'b000000011100;
		z[1488] = 3'b010;
		y[1489] = 12'b100001010111;
		z[1489] = 3'b000;
		y[1490] = 12'b001110110001;
		z[1490] = 3'b101;
		y[1491] = 12'b011010000011;
		z[1491] = 3'b110;
		y[1492] = 12'b001010101101;
		z[1492] = 3'b000;
		y[1493] = 12'b100001011100;
		z[1493] = 3'b101;
		y[1494] = 12'b100000110001;
		z[1494] = 3'b000;
		y[1495] = 12'b100101011001;
		z[1495] = 3'b110;
		y[1496] = 12'b101011100010;
		z[1496] = 3'b101;
		y[1497] = 12'b110001111001;
		z[1497] = 3'b001;
		y[1498] = 12'b000101001000;
		z[1498] = 3'b101;
		y[1499] = 12'b100101010010;
		z[1499] = 3'b011;
		y[1500] = 12'b001011011010;
		z[1500] = 3'b111;
		y[1501] = 12'b010101011010;
		z[1501] = 3'b110;
		y[1502] = 12'b010111001010;
		z[1502] = 3'b001;
		y[1503] = 12'b010101011010;
		z[1503] = 3'b100;
		y[1504] = 12'b001111111111;
		z[1504] = 3'b110;
		y[1505] = 12'b010011010111;
		z[1505] = 3'b011;
		y[1506] = 12'b100010011101;
		z[1506] = 3'b101;
		y[1507] = 12'b111010101000;
		z[1507] = 3'b010;
		y[1508] = 12'b111000110100;
		z[1508] = 3'b000;
		y[1509] = 12'b001000101001;
		z[1509] = 3'b011;
		y[1510] = 12'b110001100101;
		z[1510] = 3'b100;
		y[1511] = 12'b010110011101;
		z[1511] = 3'b001;
		y[1512] = 12'b011101111010;
		z[1512] = 3'b111;
		y[1513] = 12'b011000001001;
		z[1513] = 3'b100;
		y[1514] = 12'b110100100100;
		z[1514] = 3'b101;
		y[1515] = 12'b001011110011;
		z[1515] = 3'b010;
		y[1516] = 12'b101110111100;
		z[1516] = 3'b000;
		y[1517] = 12'b010110110110;
		z[1517] = 3'b110;
		y[1518] = 12'b001001011100;
		z[1518] = 3'b110;
		y[1519] = 12'b011100001011;
		z[1519] = 3'b000;
		y[1520] = 12'b011101101010;
		z[1520] = 3'b010;
		y[1521] = 12'b011001110110;
		z[1521] = 3'b101;
		y[1522] = 12'b100011111111;
		z[1522] = 3'b100;
		y[1523] = 12'b000101011011;
		z[1523] = 3'b110;
		y[1524] = 12'b010110111111;
		z[1524] = 3'b110;
		y[1525] = 12'b011011100101;
		z[1525] = 3'b000;
		y[1526] = 12'b000111100010;
		z[1526] = 3'b111;
		y[1527] = 12'b011110011001;
		z[1527] = 3'b010;
		y[1528] = 12'b100100101101;
		z[1528] = 3'b011;
		y[1529] = 12'b010100001111;
		z[1529] = 3'b010;
		y[1530] = 12'b000000101100;
		z[1530] = 3'b011;
		y[1531] = 12'b000000001000;
		z[1531] = 3'b101;
		y[1532] = 12'b010101011011;
		z[1532] = 3'b110;
		y[1533] = 12'b011011100001;
		z[1533] = 3'b110;
		y[1534] = 12'b001111000011;
		z[1534] = 3'b110;
		y[1535] = 12'b110100010100;
		z[1535] = 3'b000;
		y[1536] = 12'b110001110000;
		z[1536] = 3'b000;
		y[1537] = 12'b010010000100;
		z[1537] = 3'b000;
		y[1538] = 12'b001100011111;
		z[1538] = 3'b000;
		y[1539] = 12'b111011011011;
		z[1539] = 3'b000;
		y[1540] = 12'b111011111001;
		z[1540] = 3'b011;
		y[1541] = 12'b100011001000;
		z[1541] = 3'b101;
		y[1542] = 12'b110010111000;
		z[1542] = 3'b111;
		y[1543] = 12'b000010000011;
		z[1543] = 3'b000;
		y[1544] = 12'b010100001001;
		z[1544] = 3'b100;
		y[1545] = 12'b011110110010;
		z[1545] = 3'b101;
		y[1546] = 12'b000011101011;
		z[1546] = 3'b100;
		y[1547] = 12'b001111101000;
		z[1547] = 3'b010;
		y[1548] = 12'b111101010110;
		z[1548] = 3'b101;
		y[1549] = 12'b010010000111;
		z[1549] = 3'b010;
		y[1550] = 12'b110010110101;
		z[1550] = 3'b001;
		y[1551] = 12'b010110010100;
		z[1551] = 3'b111;
		y[1552] = 12'b010011111010;
		z[1552] = 3'b001;
		y[1553] = 12'b101100100010;
		z[1553] = 3'b001;
		y[1554] = 12'b101010100010;
		z[1554] = 3'b111;
		y[1555] = 12'b000101110101;
		z[1555] = 3'b011;
		y[1556] = 12'b110110011011;
		z[1556] = 3'b010;
		y[1557] = 12'b000111011101;
		z[1557] = 3'b000;
		y[1558] = 12'b001001110100;
		z[1558] = 3'b101;
		y[1559] = 12'b100111100000;
		z[1559] = 3'b011;
		y[1560] = 12'b011101111101;
		z[1560] = 3'b000;
		y[1561] = 12'b010111110101;
		z[1561] = 3'b010;
		y[1562] = 12'b000111011110;
		z[1562] = 3'b011;
		y[1563] = 12'b101111010110;
		z[1563] = 3'b111;
		y[1564] = 12'b001110011100;
		z[1564] = 3'b111;
		y[1565] = 12'b001011010001;
		z[1565] = 3'b101;
		y[1566] = 12'b010100101001;
		z[1566] = 3'b100;
		y[1567] = 12'b101100101101;
		z[1567] = 3'b000;
		y[1568] = 12'b110110110001;
		z[1568] = 3'b011;
		y[1569] = 12'b110101100011;
		z[1569] = 3'b011;
		y[1570] = 12'b100101100001;
		z[1570] = 3'b110;
		y[1571] = 12'b001011101001;
		z[1571] = 3'b000;
		y[1572] = 12'b101001011000;
		z[1572] = 3'b011;
		y[1573] = 12'b110011001101;
		z[1573] = 3'b100;
		y[1574] = 12'b110011010010;
		z[1574] = 3'b111;
		y[1575] = 12'b010111010111;
		z[1575] = 3'b010;
		y[1576] = 12'b111000100010;
		z[1576] = 3'b000;
		y[1577] = 12'b001011001101;
		z[1577] = 3'b100;
		y[1578] = 12'b011011010110;
		z[1578] = 3'b110;
		y[1579] = 12'b010000110011;
		z[1579] = 3'b100;
		y[1580] = 12'b111110001000;
		z[1580] = 3'b000;
		y[1581] = 12'b100010001100;
		z[1581] = 3'b001;
		y[1582] = 12'b100111100100;
		z[1582] = 3'b000;
		y[1583] = 12'b001000010011;
		z[1583] = 3'b001;
		y[1584] = 12'b010110101110;
		z[1584] = 3'b011;
		y[1585] = 12'b110110100011;
		z[1585] = 3'b100;
		y[1586] = 12'b010011000011;
		z[1586] = 3'b111;
		y[1587] = 12'b111001011111;
		z[1587] = 3'b011;
		y[1588] = 12'b101011001000;
		z[1588] = 3'b111;
		y[1589] = 12'b010000100000;
		z[1589] = 3'b101;
		y[1590] = 12'b100111100100;
		z[1590] = 3'b010;
		y[1591] = 12'b101101010110;
		z[1591] = 3'b111;
		y[1592] = 12'b000001000101;
		z[1592] = 3'b110;
		y[1593] = 12'b010110000001;
		z[1593] = 3'b111;
		y[1594] = 12'b000101101100;
		z[1594] = 3'b111;
		y[1595] = 12'b100100100101;
		z[1595] = 3'b001;
		y[1596] = 12'b000001111110;
		z[1596] = 3'b101;
		y[1597] = 12'b000011111101;
		z[1597] = 3'b100;
		y[1598] = 12'b110100001111;
		z[1598] = 3'b000;
		y[1599] = 12'b101010101100;
		z[1599] = 3'b010;
		y[1600] = 12'b010001001000;
		z[1600] = 3'b101;
		y[1601] = 12'b000001010100;
		z[1601] = 3'b001;
		y[1602] = 12'b101001011110;
		z[1602] = 3'b101;
		y[1603] = 12'b000001100000;
		z[1603] = 3'b001;
		y[1604] = 12'b000001001101;
		z[1604] = 3'b111;
		y[1605] = 12'b110100010110;
		z[1605] = 3'b100;
		y[1606] = 12'b001101111111;
		z[1606] = 3'b001;
		y[1607] = 12'b001001010011;
		z[1607] = 3'b000;
		y[1608] = 12'b011111010011;
		z[1608] = 3'b001;
		y[1609] = 12'b010000000110;
		z[1609] = 3'b101;
		y[1610] = 12'b111000101001;
		z[1610] = 3'b111;
		y[1611] = 12'b101010100010;
		z[1611] = 3'b111;
		y[1612] = 12'b110110011010;
		z[1612] = 3'b010;
		y[1613] = 12'b011110100111;
		z[1613] = 3'b011;
		y[1614] = 12'b001001011101;
		z[1614] = 3'b101;
		y[1615] = 12'b111101101101;
		z[1615] = 3'b000;
		y[1616] = 12'b110111010100;
		z[1616] = 3'b010;
		y[1617] = 12'b010000100000;
		z[1617] = 3'b100;
		y[1618] = 12'b100010100100;
		z[1618] = 3'b010;
		y[1619] = 12'b110110000101;
		z[1619] = 3'b011;
		y[1620] = 12'b001111001110;
		z[1620] = 3'b011;
		y[1621] = 12'b100000100101;
		z[1621] = 3'b110;
		y[1622] = 12'b100101100101;
		z[1622] = 3'b011;
		y[1623] = 12'b110010101010;
		z[1623] = 3'b010;
		y[1624] = 12'b010110011101;
		z[1624] = 3'b100;
		y[1625] = 12'b101010110011;
		z[1625] = 3'b100;
		y[1626] = 12'b100110001111;
		z[1626] = 3'b111;
		y[1627] = 12'b011101110100;
		z[1627] = 3'b111;
		y[1628] = 12'b011010100010;
		z[1628] = 3'b001;
		y[1629] = 12'b011111001011;
		z[1629] = 3'b001;
		y[1630] = 12'b010100011000;
		z[1630] = 3'b111;
		y[1631] = 12'b101101001001;
		z[1631] = 3'b101;
		y[1632] = 12'b000101110101;
		z[1632] = 3'b011;
		y[1633] = 12'b101000011010;
		z[1633] = 3'b110;
		y[1634] = 12'b111000010001;
		z[1634] = 3'b010;
		y[1635] = 12'b001001000011;
		z[1635] = 3'b101;
		y[1636] = 12'b001101010011;
		z[1636] = 3'b101;
		y[1637] = 12'b010001101010;
		z[1637] = 3'b111;
		y[1638] = 12'b010001101101;
		z[1638] = 3'b001;
		y[1639] = 12'b011000010100;
		z[1639] = 3'b100;
		y[1640] = 12'b110110110010;
		z[1640] = 3'b110;
		y[1641] = 12'b010001111101;
		z[1641] = 3'b110;
		y[1642] = 12'b011001110010;
		z[1642] = 3'b101;
		y[1643] = 12'b101010010111;
		z[1643] = 3'b000;
		y[1644] = 12'b101010111110;
		z[1644] = 3'b011;
		y[1645] = 12'b010101110110;
		z[1645] = 3'b010;
		y[1646] = 12'b011100101000;
		z[1646] = 3'b010;
		y[1647] = 12'b011111101111;
		z[1647] = 3'b001;
		y[1648] = 12'b111111101001;
		z[1648] = 3'b110;
		y[1649] = 12'b010001100100;
		z[1649] = 3'b010;
		y[1650] = 12'b101000001111;
		z[1650] = 3'b001;
		y[1651] = 12'b110000110000;
		z[1651] = 3'b100;
		y[1652] = 12'b101001110010;
		z[1652] = 3'b000;
		y[1653] = 12'b100101101110;
		z[1653] = 3'b101;
		y[1654] = 12'b111001100100;
		z[1654] = 3'b010;
		y[1655] = 12'b101110001111;
		z[1655] = 3'b000;
		y[1656] = 12'b000110110011;
		z[1656] = 3'b101;
		y[1657] = 12'b110011000001;
		z[1657] = 3'b011;
		y[1658] = 12'b001100111000;
		z[1658] = 3'b000;
		y[1659] = 12'b110001111011;
		z[1659] = 3'b001;
		y[1660] = 12'b001010001010;
		z[1660] = 3'b010;
		y[1661] = 12'b110000010011;
		z[1661] = 3'b100;
		y[1662] = 12'b110111001001;
		z[1662] = 3'b010;
		y[1663] = 12'b000100110001;
		z[1663] = 3'b110;
		y[1664] = 12'b100001000011;
		z[1664] = 3'b110;
		y[1665] = 12'b011101111100;
		z[1665] = 3'b011;
		y[1666] = 12'b110000000000;
		z[1666] = 3'b001;
		y[1667] = 12'b100110101000;
		z[1667] = 3'b110;
		y[1668] = 12'b111011100100;
		z[1668] = 3'b011;
		y[1669] = 12'b010110001111;
		z[1669] = 3'b101;
		y[1670] = 12'b010000100010;
		z[1670] = 3'b001;
		y[1671] = 12'b100000101110;
		z[1671] = 3'b110;
		y[1672] = 12'b001101000111;
		z[1672] = 3'b011;
		y[1673] = 12'b100111011000;
		z[1673] = 3'b111;
		y[1674] = 12'b010010000000;
		z[1674] = 3'b101;
		y[1675] = 12'b110010111010;
		z[1675] = 3'b101;
		y[1676] = 12'b000110101000;
		z[1676] = 3'b001;
		y[1677] = 12'b001111111000;
		z[1677] = 3'b111;
		y[1678] = 12'b001000100110;
		z[1678] = 3'b101;
		y[1679] = 12'b110000100001;
		z[1679] = 3'b101;
		y[1680] = 12'b101000101101;
		z[1680] = 3'b011;
		y[1681] = 12'b000101101100;
		z[1681] = 3'b111;
		y[1682] = 12'b110011101000;
		z[1682] = 3'b110;
		y[1683] = 12'b000000011110;
		z[1683] = 3'b011;
		y[1684] = 12'b111101101111;
		z[1684] = 3'b000;
		y[1685] = 12'b100010100101;
		z[1685] = 3'b000;
		y[1686] = 12'b011111111011;
		z[1686] = 3'b011;
		y[1687] = 12'b100100100100;
		z[1687] = 3'b000;
		y[1688] = 12'b010110010011;
		z[1688] = 3'b111;
		y[1689] = 12'b111111101000;
		z[1689] = 3'b101;
		y[1690] = 12'b110101001111;
		z[1690] = 3'b011;
		y[1691] = 12'b001000111010;
		z[1691] = 3'b110;
		y[1692] = 12'b011110110010;
		z[1692] = 3'b110;
		y[1693] = 12'b111100000011;
		z[1693] = 3'b000;
		y[1694] = 12'b111000010110;
		z[1694] = 3'b111;
		y[1695] = 12'b101101010011;
		z[1695] = 3'b001;
		y[1696] = 12'b100100000001;
		z[1696] = 3'b010;
		y[1697] = 12'b110011010000;
		z[1697] = 3'b110;
		y[1698] = 12'b000001101010;
		z[1698] = 3'b011;
		y[1699] = 12'b001101100011;
		z[1699] = 3'b000;
		y[1700] = 12'b101010111010;
		z[1700] = 3'b101;
		y[1701] = 12'b011111010100;
		z[1701] = 3'b100;
		y[1702] = 12'b110001010101;
		z[1702] = 3'b101;
		y[1703] = 12'b100100111111;
		z[1703] = 3'b001;
		y[1704] = 12'b100001011100;
		z[1704] = 3'b001;
		y[1705] = 12'b001101001001;
		z[1705] = 3'b000;
		y[1706] = 12'b100011011011;
		z[1706] = 3'b011;
		y[1707] = 12'b010111000100;
		z[1707] = 3'b001;
		y[1708] = 12'b010101001011;
		z[1708] = 3'b011;
		y[1709] = 12'b110010010110;
		z[1709] = 3'b000;
		y[1710] = 12'b011001111001;
		z[1710] = 3'b110;
		y[1711] = 12'b100000111011;
		z[1711] = 3'b011;
		y[1712] = 12'b010001100000;
		z[1712] = 3'b100;
		y[1713] = 12'b110001110010;
		z[1713] = 3'b110;
		y[1714] = 12'b011000000100;
		z[1714] = 3'b011;
		y[1715] = 12'b110001000010;
		z[1715] = 3'b010;
		y[1716] = 12'b011011111001;
		z[1716] = 3'b010;
		y[1717] = 12'b010111010011;
		z[1717] = 3'b010;
		y[1718] = 12'b011010101110;
		z[1718] = 3'b100;
		y[1719] = 12'b110100001101;
		z[1719] = 3'b001;
		y[1720] = 12'b110101101000;
		z[1720] = 3'b001;
		y[1721] = 12'b001000111011;
		z[1721] = 3'b010;
		y[1722] = 12'b100011100010;
		z[1722] = 3'b011;
		y[1723] = 12'b111010010001;
		z[1723] = 3'b011;
		y[1724] = 12'b111000110110;
		z[1724] = 3'b100;
		y[1725] = 12'b010000000011;
		z[1725] = 3'b010;
		y[1726] = 12'b100001011001;
		z[1726] = 3'b011;
		y[1727] = 12'b100001100010;
		z[1727] = 3'b011;
		y[1728] = 12'b010010111100;
		z[1728] = 3'b100;
		y[1729] = 12'b101100011010;
		z[1729] = 3'b100;
		y[1730] = 12'b100101110101;
		z[1730] = 3'b000;
		y[1731] = 12'b110011000001;
		z[1731] = 3'b001;
		y[1732] = 12'b100100100000;
		z[1732] = 3'b111;
		y[1733] = 12'b000010001100;
		z[1733] = 3'b011;
		y[1734] = 12'b000001011000;
		z[1734] = 3'b011;
		y[1735] = 12'b101011101000;
		z[1735] = 3'b110;
		y[1736] = 12'b011111011001;
		z[1736] = 3'b001;
		y[1737] = 12'b010111100010;
		z[1737] = 3'b100;
		y[1738] = 12'b111000110111;
		z[1738] = 3'b100;
		y[1739] = 12'b110101001010;
		z[1739] = 3'b011;
		y[1740] = 12'b011101101100;
		z[1740] = 3'b111;
		y[1741] = 12'b010000010001;
		z[1741] = 3'b010;
		y[1742] = 12'b110110110110;
		z[1742] = 3'b111;
		y[1743] = 12'b010000100101;
		z[1743] = 3'b110;
		y[1744] = 12'b010011010101;
		z[1744] = 3'b111;
		y[1745] = 12'b100000011000;
		z[1745] = 3'b011;
		y[1746] = 12'b000100010100;
		z[1746] = 3'b011;
		y[1747] = 12'b011101011001;
		z[1747] = 3'b110;
		y[1748] = 12'b101000011010;
		z[1748] = 3'b000;
		y[1749] = 12'b101001110001;
		z[1749] = 3'b000;
		y[1750] = 12'b001110001011;
		z[1750] = 3'b010;
		y[1751] = 12'b001010001101;
		z[1751] = 3'b010;
		y[1752] = 12'b100111000111;
		z[1752] = 3'b011;
		y[1753] = 12'b011101111110;
		z[1753] = 3'b000;
		y[1754] = 12'b110010001010;
		z[1754] = 3'b110;
		y[1755] = 12'b000110001010;
		z[1755] = 3'b011;
		y[1756] = 12'b011110011010;
		z[1756] = 3'b100;
		y[1757] = 12'b100010100000;
		z[1757] = 3'b110;
		y[1758] = 12'b110110001101;
		z[1758] = 3'b101;
		y[1759] = 12'b011001001011;
		z[1759] = 3'b100;
		y[1760] = 12'b100100110001;
		z[1760] = 3'b010;
		y[1761] = 12'b101000101111;
		z[1761] = 3'b101;
		y[1762] = 12'b001010001111;
		z[1762] = 3'b010;
		y[1763] = 12'b110001101001;
		z[1763] = 3'b011;
		y[1764] = 12'b111100110110;
		z[1764] = 3'b010;
		y[1765] = 12'b011010100111;
		z[1765] = 3'b101;
		y[1766] = 12'b111010111010;
		z[1766] = 3'b000;
		y[1767] = 12'b011010111000;
		z[1767] = 3'b111;
		y[1768] = 12'b011010100010;
		z[1768] = 3'b011;
		y[1769] = 12'b101011110100;
		z[1769] = 3'b110;
		y[1770] = 12'b101000001111;
		z[1770] = 3'b110;
		y[1771] = 12'b101110000100;
		z[1771] = 3'b011;
		y[1772] = 12'b011110000010;
		z[1772] = 3'b010;
		y[1773] = 12'b111001011011;
		z[1773] = 3'b010;
		y[1774] = 12'b100110000010;
		z[1774] = 3'b001;
		y[1775] = 12'b110110101000;
		z[1775] = 3'b100;
		y[1776] = 12'b101111001000;
		z[1776] = 3'b111;
		y[1777] = 12'b000101010101;
		z[1777] = 3'b111;
		y[1778] = 12'b011010111010;
		z[1778] = 3'b111;
		y[1779] = 12'b110010010110;
		z[1779] = 3'b001;
		y[1780] = 12'b111010101110;
		z[1780] = 3'b010;
		y[1781] = 12'b111000011011;
		z[1781] = 3'b101;
		y[1782] = 12'b000101011100;
		z[1782] = 3'b110;
		y[1783] = 12'b100001110111;
		z[1783] = 3'b100;
		y[1784] = 12'b000111010101;
		z[1784] = 3'b000;
		y[1785] = 12'b000100111100;
		z[1785] = 3'b001;
		y[1786] = 12'b100000011001;
		z[1786] = 3'b110;
		y[1787] = 12'b111111110111;
		z[1787] = 3'b011;
		y[1788] = 12'b111111011010;
		z[1788] = 3'b111;
		y[1789] = 12'b100000001011;
		z[1789] = 3'b110;
		y[1790] = 12'b101110111011;
		z[1790] = 3'b011;
		y[1791] = 12'b111000110110;
		z[1791] = 3'b101;
		y[1792] = 12'b000011010010;
		z[1792] = 3'b010;
		y[1793] = 12'b010111011001;
		z[1793] = 3'b110;
		y[1794] = 12'b001110010000;
		z[1794] = 3'b001;
		y[1795] = 12'b110101100110;
		z[1795] = 3'b100;
		y[1796] = 12'b001000000101;
		z[1796] = 3'b100;
		y[1797] = 12'b111001000100;
		z[1797] = 3'b100;
		y[1798] = 12'b000010011101;
		z[1798] = 3'b010;
		y[1799] = 12'b111000100011;
		z[1799] = 3'b000;
		y[1800] = 12'b100100011101;
		z[1800] = 3'b011;
		y[1801] = 12'b000000011011;
		z[1801] = 3'b111;
		y[1802] = 12'b110001001110;
		z[1802] = 3'b110;
		y[1803] = 12'b101101110111;
		z[1803] = 3'b100;
		y[1804] = 12'b100100011111;
		z[1804] = 3'b110;
		y[1805] = 12'b101100110101;
		z[1805] = 3'b100;
		y[1806] = 12'b100010111100;
		z[1806] = 3'b011;
		y[1807] = 12'b101111111111;
		z[1807] = 3'b111;
		y[1808] = 12'b101110001110;
		z[1808] = 3'b100;
		y[1809] = 12'b000010010010;
		z[1809] = 3'b011;
		y[1810] = 12'b101101111100;
		z[1810] = 3'b111;
		y[1811] = 12'b110010100111;
		z[1811] = 3'b000;
		y[1812] = 12'b000000010101;
		z[1812] = 3'b110;
		y[1813] = 12'b111100101100;
		z[1813] = 3'b100;
		y[1814] = 12'b111101100110;
		z[1814] = 3'b000;
		y[1815] = 12'b000000010010;
		z[1815] = 3'b000;
		y[1816] = 12'b010001001001;
		z[1816] = 3'b000;
		y[1817] = 12'b001111110000;
		z[1817] = 3'b110;
		y[1818] = 12'b010011110111;
		z[1818] = 3'b100;
		y[1819] = 12'b011000110111;
		z[1819] = 3'b010;
		y[1820] = 12'b011111011001;
		z[1820] = 3'b011;
		y[1821] = 12'b011101001111;
		z[1821] = 3'b111;
		y[1822] = 12'b001011011001;
		z[1822] = 3'b011;
		y[1823] = 12'b000111110001;
		z[1823] = 3'b000;
		y[1824] = 12'b110010100100;
		z[1824] = 3'b101;
		y[1825] = 12'b001101001111;
		z[1825] = 3'b000;
		y[1826] = 12'b010001111100;
		z[1826] = 3'b100;
		y[1827] = 12'b101011000111;
		z[1827] = 3'b011;
		y[1828] = 12'b010101001101;
		z[1828] = 3'b000;
		y[1829] = 12'b000101010011;
		z[1829] = 3'b110;
		y[1830] = 12'b011101111010;
		z[1830] = 3'b001;
		y[1831] = 12'b000000101101;
		z[1831] = 3'b101;
		y[1832] = 12'b000011110011;
		z[1832] = 3'b000;
		y[1833] = 12'b100000100001;
		z[1833] = 3'b000;
		y[1834] = 12'b110000101001;
		z[1834] = 3'b001;
		y[1835] = 12'b110111101010;
		z[1835] = 3'b010;
		y[1836] = 12'b010011010000;
		z[1836] = 3'b010;
		y[1837] = 12'b100011100111;
		z[1837] = 3'b001;
		y[1838] = 12'b111100011000;
		z[1838] = 3'b110;
		y[1839] = 12'b010101000011;
		z[1839] = 3'b100;
		y[1840] = 12'b010111001100;
		z[1840] = 3'b011;
		y[1841] = 12'b000100111000;
		z[1841] = 3'b010;
		y[1842] = 12'b000010001110;
		z[1842] = 3'b100;
		y[1843] = 12'b101001010100;
		z[1843] = 3'b001;
		y[1844] = 12'b110110101000;
		z[1844] = 3'b011;
		y[1845] = 12'b011011010001;
		z[1845] = 3'b010;
		y[1846] = 12'b010111001000;
		z[1846] = 3'b100;
		y[1847] = 12'b001110100101;
		z[1847] = 3'b000;
		y[1848] = 12'b010001110010;
		z[1848] = 3'b011;
		y[1849] = 12'b110101100101;
		z[1849] = 3'b011;
		y[1850] = 12'b101011011100;
		z[1850] = 3'b001;
		y[1851] = 12'b011000101100;
		z[1851] = 3'b110;
		y[1852] = 12'b110101100110;
		z[1852] = 3'b011;
		y[1853] = 12'b001100000100;
		z[1853] = 3'b111;
		y[1854] = 12'b101010110110;
		z[1854] = 3'b111;
		y[1855] = 12'b110010001111;
		z[1855] = 3'b101;
		y[1856] = 12'b110110001011;
		z[1856] = 3'b001;
		y[1857] = 12'b110101001001;
		z[1857] = 3'b100;
		y[1858] = 12'b000011100111;
		z[1858] = 3'b101;
		y[1859] = 12'b001110101011;
		z[1859] = 3'b101;
		y[1860] = 12'b101010100100;
		z[1860] = 3'b011;
		y[1861] = 12'b111111000100;
		z[1861] = 3'b010;
		y[1862] = 12'b100100010000;
		z[1862] = 3'b011;
		y[1863] = 12'b000110000101;
		z[1863] = 3'b101;
		y[1864] = 12'b001101110010;
		z[1864] = 3'b110;
		y[1865] = 12'b010111111001;
		z[1865] = 3'b010;
		y[1866] = 12'b011110111101;
		z[1866] = 3'b001;
		y[1867] = 12'b010000011111;
		z[1867] = 3'b111;
		y[1868] = 12'b000000011000;
		z[1868] = 3'b001;
		y[1869] = 12'b000110110101;
		z[1869] = 3'b011;
		y[1870] = 12'b010100111100;
		z[1870] = 3'b100;
		y[1871] = 12'b001101100010;
		z[1871] = 3'b001;
		y[1872] = 12'b110001010000;
		z[1872] = 3'b010;
		y[1873] = 12'b111010111010;
		z[1873] = 3'b001;
		y[1874] = 12'b000000110100;
		z[1874] = 3'b100;
		y[1875] = 12'b010111010111;
		z[1875] = 3'b001;
		y[1876] = 12'b000001101111;
		z[1876] = 3'b100;
		y[1877] = 12'b011111000000;
		z[1877] = 3'b100;
		y[1878] = 12'b000010010000;
		z[1878] = 3'b000;
		y[1879] = 12'b110010011101;
		z[1879] = 3'b111;
		y[1880] = 12'b101101000101;
		z[1880] = 3'b111;
		y[1881] = 12'b110110110010;
		z[1881] = 3'b010;
		y[1882] = 12'b001001011010;
		z[1882] = 3'b111;
		y[1883] = 12'b101111111010;
		z[1883] = 3'b001;
		y[1884] = 12'b101100010011;
		z[1884] = 3'b110;
		y[1885] = 12'b101000011000;
		z[1885] = 3'b011;
		y[1886] = 12'b111110011011;
		z[1886] = 3'b011;
		y[1887] = 12'b010111000101;
		z[1887] = 3'b101;
		y[1888] = 12'b000101100011;
		z[1888] = 3'b111;
		y[1889] = 12'b101000001001;
		z[1889] = 3'b000;
		y[1890] = 12'b000101111110;
		z[1890] = 3'b101;
		y[1891] = 12'b110011101011;
		z[1891] = 3'b010;
		y[1892] = 12'b111111101111;
		z[1892] = 3'b010;
		y[1893] = 12'b011001001011;
		z[1893] = 3'b000;
		y[1894] = 12'b010011000101;
		z[1894] = 3'b001;
		y[1895] = 12'b011111101101;
		z[1895] = 3'b011;
		y[1896] = 12'b010100000000;
		z[1896] = 3'b011;
		y[1897] = 12'b111101011000;
		z[1897] = 3'b101;
		y[1898] = 12'b010000000001;
		z[1898] = 3'b011;
		y[1899] = 12'b100100001100;
		z[1899] = 3'b010;
		y[1900] = 12'b100100000011;
		z[1900] = 3'b000;
		y[1901] = 12'b100111001101;
		z[1901] = 3'b000;
		y[1902] = 12'b111001110111;
		z[1902] = 3'b001;
		y[1903] = 12'b010011100110;
		z[1903] = 3'b110;
		y[1904] = 12'b111000010001;
		z[1904] = 3'b111;
		y[1905] = 12'b111000111101;
		z[1905] = 3'b111;
		y[1906] = 12'b100000011100;
		z[1906] = 3'b110;
		y[1907] = 12'b101001011111;
		z[1907] = 3'b001;
		y[1908] = 12'b101010011110;
		z[1908] = 3'b110;
		y[1909] = 12'b011001010101;
		z[1909] = 3'b110;
		y[1910] = 12'b110000000101;
		z[1910] = 3'b000;
		y[1911] = 12'b010101100000;
		z[1911] = 3'b000;
		y[1912] = 12'b111110000010;
		z[1912] = 3'b101;
		y[1913] = 12'b100111101101;
		z[1913] = 3'b111;
		y[1914] = 12'b000101010001;
		z[1914] = 3'b100;
		y[1915] = 12'b111010101000;
		z[1915] = 3'b010;
		y[1916] = 12'b111111000000;
		z[1916] = 3'b011;
		y[1917] = 12'b100010001101;
		z[1917] = 3'b010;
		y[1918] = 12'b001010100000;
		z[1918] = 3'b000;
		y[1919] = 12'b111011010001;
		z[1919] = 3'b001;
		y[1920] = 12'b001111111100;
		z[1920] = 3'b111;
		y[1921] = 12'b100111010110;
		z[1921] = 3'b111;
		y[1922] = 12'b111011011011;
		z[1922] = 3'b011;
		y[1923] = 12'b111000110001;
		z[1923] = 3'b100;
		y[1924] = 12'b110111100010;
		z[1924] = 3'b000;
		y[1925] = 12'b111011001111;
		z[1925] = 3'b000;
		y[1926] = 12'b111101010110;
		z[1926] = 3'b000;
		y[1927] = 12'b110110000111;
		z[1927] = 3'b100;
		y[1928] = 12'b100001110110;
		z[1928] = 3'b010;
		y[1929] = 12'b100100011100;
		z[1929] = 3'b101;
		y[1930] = 12'b100110010110;
		z[1930] = 3'b110;
		y[1931] = 12'b010010010111;
		z[1931] = 3'b100;
		y[1932] = 12'b000011010110;
		z[1932] = 3'b101;
		y[1933] = 12'b001000010111;
		z[1933] = 3'b011;
		y[1934] = 12'b111011100010;
		z[1934] = 3'b001;
		y[1935] = 12'b001100101011;
		z[1935] = 3'b010;
		y[1936] = 12'b000010011010;
		z[1936] = 3'b000;
		y[1937] = 12'b101010001110;
		z[1937] = 3'b011;
		y[1938] = 12'b010010110001;
		z[1938] = 3'b001;
		y[1939] = 12'b001100011110;
		z[1939] = 3'b010;
		y[1940] = 12'b101100001011;
		z[1940] = 3'b011;
		y[1941] = 12'b110010001100;
		z[1941] = 3'b010;
		y[1942] = 12'b100110011011;
		z[1942] = 3'b000;
		y[1943] = 12'b000110000011;
		z[1943] = 3'b001;
		y[1944] = 12'b110010110011;
		z[1944] = 3'b010;
		y[1945] = 12'b100010010110;
		z[1945] = 3'b010;
		y[1946] = 12'b000110001110;
		z[1946] = 3'b001;
		y[1947] = 12'b110101110011;
		z[1947] = 3'b011;
		y[1948] = 12'b000001010110;
		z[1948] = 3'b010;
		y[1949] = 12'b100101111110;
		z[1949] = 3'b011;
		y[1950] = 12'b100001110010;
		z[1950] = 3'b001;
		y[1951] = 12'b000111011001;
		z[1951] = 3'b111;
		y[1952] = 12'b111010100101;
		z[1952] = 3'b000;
		y[1953] = 12'b110011000101;
		z[1953] = 3'b111;
		y[1954] = 12'b010001111010;
		z[1954] = 3'b010;
		y[1955] = 12'b001100111001;
		z[1955] = 3'b000;
		y[1956] = 12'b100001000001;
		z[1956] = 3'b001;
		y[1957] = 12'b110011100101;
		z[1957] = 3'b000;
		y[1958] = 12'b101011110100;
		z[1958] = 3'b111;
		y[1959] = 12'b110001010100;
		z[1959] = 3'b111;
		y[1960] = 12'b000010000110;
		z[1960] = 3'b001;
		y[1961] = 12'b000110000110;
		z[1961] = 3'b111;
		y[1962] = 12'b100100100101;
		z[1962] = 3'b000;
		y[1963] = 12'b110110011000;
		z[1963] = 3'b001;
		y[1964] = 12'b000000110000;
		z[1964] = 3'b010;
		y[1965] = 12'b110001001110;
		z[1965] = 3'b100;
		y[1966] = 12'b100010001110;
		z[1966] = 3'b101;
		y[1967] = 12'b101101100100;
		z[1967] = 3'b010;
		y[1968] = 12'b000000001100;
		z[1968] = 3'b000;
		y[1969] = 12'b011010010010;
		z[1969] = 3'b011;
		y[1970] = 12'b000001000010;
		z[1970] = 3'b000;
		y[1971] = 12'b100010011101;
		z[1971] = 3'b101;
		y[1972] = 12'b010101011000;
		z[1972] = 3'b010;
		y[1973] = 12'b000101101000;
		z[1973] = 3'b010;
		y[1974] = 12'b100101010100;
		z[1974] = 3'b010;
		y[1975] = 12'b011100011100;
		z[1975] = 3'b001;
		y[1976] = 12'b010101111110;
		z[1976] = 3'b111;
		y[1977] = 12'b111001000101;
		z[1977] = 3'b111;
		y[1978] = 12'b010110001111;
		z[1978] = 3'b100;
		y[1979] = 12'b110000001001;
		z[1979] = 3'b111;
		y[1980] = 12'b110011111001;
		z[1980] = 3'b100;
		y[1981] = 12'b000001011001;
		z[1981] = 3'b010;
		y[1982] = 12'b101001110010;
		z[1982] = 3'b101;
		y[1983] = 12'b110000100010;
		z[1983] = 3'b001;
		y[1984] = 12'b111000110001;
		z[1984] = 3'b010;
		y[1985] = 12'b000101000101;
		z[1985] = 3'b100;
		y[1986] = 12'b010111001111;
		z[1986] = 3'b101;
		y[1987] = 12'b010010011101;
		z[1987] = 3'b010;
		y[1988] = 12'b101000011010;
		z[1988] = 3'b101;
		y[1989] = 12'b010001000111;
		z[1989] = 3'b100;
		y[1990] = 12'b101111011100;
		z[1990] = 3'b111;
		y[1991] = 12'b111010101011;
		z[1991] = 3'b111;
		y[1992] = 12'b111101111010;
		z[1992] = 3'b000;
		y[1993] = 12'b001010111111;
		z[1993] = 3'b011;
		y[1994] = 12'b011111101011;
		z[1994] = 3'b101;
		y[1995] = 12'b011110001111;
		z[1995] = 3'b011;
		y[1996] = 12'b011101000101;
		z[1996] = 3'b100;
		y[1997] = 12'b100000100000;
		z[1997] = 3'b100;
		y[1998] = 12'b010111111100;
		z[1998] = 3'b000;
		y[1999] = 12'b101110101110;
		z[1999] = 3'b111;
		y[2000] = 12'b011000110111;
		z[2000] = 3'b100;
		y[2001] = 12'b100010010110;
		z[2001] = 3'b001;
		y[2002] = 12'b110100000010;
		z[2002] = 3'b101;
		y[2003] = 12'b100110110101;
		z[2003] = 3'b010;
		y[2004] = 12'b000010001011;
		z[2004] = 3'b011;
		y[2005] = 12'b010000011110;
		z[2005] = 3'b001;
		y[2006] = 12'b010111011111;
		z[2006] = 3'b000;
		y[2007] = 12'b000100010111;
		z[2007] = 3'b000;
		y[2008] = 12'b100000000111;
		z[2008] = 3'b001;
		y[2009] = 12'b110000110101;
		z[2009] = 3'b000;
		y[2010] = 12'b100111100011;
		z[2010] = 3'b111;
		y[2011] = 12'b001010101110;
		z[2011] = 3'b111;
		y[2012] = 12'b101101101000;
		z[2012] = 3'b000;
		y[2013] = 12'b000001111110;
		z[2013] = 3'b111;
		y[2014] = 12'b000101001111;
		z[2014] = 3'b000;
		y[2015] = 12'b101110111000;
		z[2015] = 3'b101;
		y[2016] = 12'b010101110011;
		z[2016] = 3'b110;
		y[2017] = 12'b000110101111;
		z[2017] = 3'b101;
		y[2018] = 12'b111000101010;
		z[2018] = 3'b100;
		y[2019] = 12'b101101100100;
		z[2019] = 3'b110;
		y[2020] = 12'b110101111101;
		z[2020] = 3'b000;
		y[2021] = 12'b110100010111;
		z[2021] = 3'b110;
		y[2022] = 12'b110000001110;
		z[2022] = 3'b010;
		y[2023] = 12'b000110001111;
		z[2023] = 3'b110;
		y[2024] = 12'b100000000010;
		z[2024] = 3'b001;
		y[2025] = 12'b110100000100;
		z[2025] = 3'b101;
		y[2026] = 12'b100111011100;
		z[2026] = 3'b010;
		y[2027] = 12'b010011100011;
		z[2027] = 3'b101;
		y[2028] = 12'b111010010011;
		z[2028] = 3'b101;
		y[2029] = 12'b100110100000;
		z[2029] = 3'b100;
		y[2030] = 12'b001101100010;
		z[2030] = 3'b011;
		y[2031] = 12'b100001011001;
		z[2031] = 3'b100;
		y[2032] = 12'b111011101010;
		z[2032] = 3'b000;
		y[2033] = 12'b110001010000;
		z[2033] = 3'b110;
		y[2034] = 12'b111000000100;
		z[2034] = 3'b010;
		y[2035] = 12'b011000101011;
		z[2035] = 3'b001;
		y[2036] = 12'b111001001101;
		z[2036] = 3'b111;
		y[2037] = 12'b011100001111;
		z[2037] = 3'b000;
		y[2038] = 12'b011010010011;
		z[2038] = 3'b100;
		y[2039] = 12'b111011010101;
		z[2039] = 3'b011;
		y[2040] = 12'b001110011100;
		z[2040] = 3'b101;
		y[2041] = 12'b110110100011;
		z[2041] = 3'b001;
		y[2042] = 12'b111111001101;
		z[2042] = 3'b100;
		y[2043] = 12'b111110010111;
		z[2043] = 3'b101;
		y[2044] = 12'b111100101111;
		z[2044] = 3'b101;
		y[2045] = 12'b010010111101;
		z[2045] = 3'b111;
		y[2046] = 12'b100101110010;
		z[2046] = 3'b111;
		y[2047] = 12'b100010000000;
		z[2047] = 3'b100;
		y[2048] = 12'b000100100101;
		z[2048] = 3'b100;
		y[2049] = 12'b100110010011;
		z[2049] = 3'b101;
		y[2050] = 12'b001011111111;
		z[2050] = 3'b001;
		y[2051] = 12'b101001000100;
		z[2051] = 3'b111;
		y[2052] = 12'b100011101011;
		z[2052] = 3'b000;
		y[2053] = 12'b100101000101;
		z[2053] = 3'b111;
		y[2054] = 12'b011011000110;
		z[2054] = 3'b011;
		y[2055] = 12'b010100000001;
		z[2055] = 3'b111;
		y[2056] = 12'b111101011101;
		z[2056] = 3'b011;
		y[2057] = 12'b101100001010;
		z[2057] = 3'b110;
		y[2058] = 12'b000101101111;
		z[2058] = 3'b001;
		y[2059] = 12'b110011011100;
		z[2059] = 3'b100;
		y[2060] = 12'b100010101001;
		z[2060] = 3'b101;
		y[2061] = 12'b100110110111;
		z[2061] = 3'b111;
		y[2062] = 12'b011000111110;
		z[2062] = 3'b000;
		y[2063] = 12'b111111101001;
		z[2063] = 3'b001;
		y[2064] = 12'b110100000010;
		z[2064] = 3'b001;
		y[2065] = 12'b000001100100;
		z[2065] = 3'b101;
		y[2066] = 12'b001101100001;
		z[2066] = 3'b010;
		y[2067] = 12'b100110100000;
		z[2067] = 3'b001;
		y[2068] = 12'b111000100111;
		z[2068] = 3'b111;
		y[2069] = 12'b110000111111;
		z[2069] = 3'b011;
		y[2070] = 12'b111111111011;
		z[2070] = 3'b101;
		y[2071] = 12'b000110100101;
		z[2071] = 3'b001;
		y[2072] = 12'b111000101001;
		z[2072] = 3'b001;
		y[2073] = 12'b101011000100;
		z[2073] = 3'b000;
		y[2074] = 12'b100111101011;
		z[2074] = 3'b010;
		y[2075] = 12'b000100110101;
		z[2075] = 3'b110;
		y[2076] = 12'b101010000111;
		z[2076] = 3'b011;
		y[2077] = 12'b001100110101;
		z[2077] = 3'b110;
		y[2078] = 12'b010000000100;
		z[2078] = 3'b000;
		y[2079] = 12'b000110000101;
		z[2079] = 3'b100;
		y[2080] = 12'b110001011010;
		z[2080] = 3'b000;
		y[2081] = 12'b011000111100;
		z[2081] = 3'b011;
		y[2082] = 12'b001011101100;
		z[2082] = 3'b100;
		y[2083] = 12'b010010100100;
		z[2083] = 3'b011;
		y[2084] = 12'b010101010101;
		z[2084] = 3'b000;
		y[2085] = 12'b111101100000;
		z[2085] = 3'b001;
		y[2086] = 12'b111100010101;
		z[2086] = 3'b000;
		y[2087] = 12'b010010011101;
		z[2087] = 3'b100;
		y[2088] = 12'b111011000011;
		z[2088] = 3'b010;
		y[2089] = 12'b110111101001;
		z[2089] = 3'b000;
		y[2090] = 12'b000011110010;
		z[2090] = 3'b000;
		y[2091] = 12'b110010001011;
		z[2091] = 3'b011;
		y[2092] = 12'b110101100100;
		z[2092] = 3'b100;
		y[2093] = 12'b011001000100;
		z[2093] = 3'b010;
		y[2094] = 12'b000011000101;
		z[2094] = 3'b011;
		y[2095] = 12'b111010111101;
		z[2095] = 3'b011;
		y[2096] = 12'b100001010110;
		z[2096] = 3'b111;
		y[2097] = 12'b111011011000;
		z[2097] = 3'b110;
		y[2098] = 12'b011000101100;
		z[2098] = 3'b111;
		y[2099] = 12'b000101100111;
		z[2099] = 3'b010;
		y[2100] = 12'b111001111111;
		z[2100] = 3'b001;
		y[2101] = 12'b011110011111;
		z[2101] = 3'b110;
		y[2102] = 12'b111001101101;
		z[2102] = 3'b101;
		y[2103] = 12'b010110011101;
		z[2103] = 3'b011;
		y[2104] = 12'b000100110101;
		z[2104] = 3'b010;
		y[2105] = 12'b110011111011;
		z[2105] = 3'b110;
		y[2106] = 12'b110111100010;
		z[2106] = 3'b111;
		y[2107] = 12'b101010010010;
		z[2107] = 3'b111;
		y[2108] = 12'b010101000110;
		z[2108] = 3'b001;
		y[2109] = 12'b010011001101;
		z[2109] = 3'b001;
		y[2110] = 12'b011111000111;
		z[2110] = 3'b110;
		y[2111] = 12'b110100100111;
		z[2111] = 3'b100;
		y[2112] = 12'b001000010100;
		z[2112] = 3'b111;
		y[2113] = 12'b000101110001;
		z[2113] = 3'b100;
		y[2114] = 12'b010110011110;
		z[2114] = 3'b100;
		y[2115] = 12'b001000110100;
		z[2115] = 3'b101;
		y[2116] = 12'b110111111010;
		z[2116] = 3'b011;
		y[2117] = 12'b111110011101;
		z[2117] = 3'b100;
		y[2118] = 12'b011000010000;
		z[2118] = 3'b011;
		y[2119] = 12'b101000000000;
		z[2119] = 3'b111;
		y[2120] = 12'b111001011100;
		z[2120] = 3'b100;
		y[2121] = 12'b101001000011;
		z[2121] = 3'b111;
		y[2122] = 12'b001000110100;
		z[2122] = 3'b011;
		y[2123] = 12'b011111110100;
		z[2123] = 3'b110;
		y[2124] = 12'b001000110100;
		z[2124] = 3'b101;
		y[2125] = 12'b110111010110;
		z[2125] = 3'b011;
		y[2126] = 12'b010100000001;
		z[2126] = 3'b001;
		y[2127] = 12'b011000111110;
		z[2127] = 3'b001;
		y[2128] = 12'b000011010011;
		z[2128] = 3'b110;
		y[2129] = 12'b011100100011;
		z[2129] = 3'b010;
		y[2130] = 12'b111100101010;
		z[2130] = 3'b101;
		y[2131] = 12'b110000001110;
		z[2131] = 3'b010;
		y[2132] = 12'b001101010100;
		z[2132] = 3'b100;
		y[2133] = 12'b011110101010;
		z[2133] = 3'b010;
		y[2134] = 12'b101101001000;
		z[2134] = 3'b011;
		y[2135] = 12'b110110101000;
		z[2135] = 3'b110;
		y[2136] = 12'b110110100010;
		z[2136] = 3'b000;
		y[2137] = 12'b001010010001;
		z[2137] = 3'b010;
		y[2138] = 12'b000110111100;
		z[2138] = 3'b110;
		y[2139] = 12'b000101111010;
		z[2139] = 3'b011;
		y[2140] = 12'b101000110110;
		z[2140] = 3'b101;
		y[2141] = 12'b110110100001;
		z[2141] = 3'b000;
		y[2142] = 12'b101111100111;
		z[2142] = 3'b000;
		y[2143] = 12'b011110011001;
		z[2143] = 3'b111;
		y[2144] = 12'b101001000001;
		z[2144] = 3'b111;
		y[2145] = 12'b101111111000;
		z[2145] = 3'b101;
		y[2146] = 12'b000100001110;
		z[2146] = 3'b110;
		y[2147] = 12'b011101111010;
		z[2147] = 3'b000;
		y[2148] = 12'b011100111111;
		z[2148] = 3'b011;
		y[2149] = 12'b000110010000;
		z[2149] = 3'b111;
		y[2150] = 12'b111100110110;
		z[2150] = 3'b011;
		y[2151] = 12'b000010001010;
		z[2151] = 3'b100;
		y[2152] = 12'b011001000001;
		z[2152] = 3'b110;
		y[2153] = 12'b111110011010;
		z[2153] = 3'b000;
		y[2154] = 12'b011111111100;
		z[2154] = 3'b111;
		y[2155] = 12'b101001011000;
		z[2155] = 3'b110;
		y[2156] = 12'b000100010100;
		z[2156] = 3'b111;
		y[2157] = 12'b010110100111;
		z[2157] = 3'b001;
		y[2158] = 12'b110100011000;
		z[2158] = 3'b001;
		y[2159] = 12'b100110111100;
		z[2159] = 3'b000;
		y[2160] = 12'b101010110100;
		z[2160] = 3'b111;
		y[2161] = 12'b010100111110;
		z[2161] = 3'b101;
		y[2162] = 12'b011101010011;
		z[2162] = 3'b111;
		y[2163] = 12'b111100011110;
		z[2163] = 3'b010;
		y[2164] = 12'b111110001010;
		z[2164] = 3'b111;
		y[2165] = 12'b101100100111;
		z[2165] = 3'b000;
		y[2166] = 12'b001001101010;
		z[2166] = 3'b111;
		y[2167] = 12'b001001000100;
		z[2167] = 3'b111;
		y[2168] = 12'b111100111000;
		z[2168] = 3'b001;
		y[2169] = 12'b010010110001;
		z[2169] = 3'b001;
		y[2170] = 12'b100101111011;
		z[2170] = 3'b110;
		y[2171] = 12'b101011001110;
		z[2171] = 3'b110;
		y[2172] = 12'b001111011011;
		z[2172] = 3'b000;
		y[2173] = 12'b000111001101;
		z[2173] = 3'b110;
		y[2174] = 12'b001101100001;
		z[2174] = 3'b100;
		y[2175] = 12'b001110010010;
		z[2175] = 3'b111;
		y[2176] = 12'b001100000101;
		z[2176] = 3'b000;
		y[2177] = 12'b011000110011;
		z[2177] = 3'b100;
		y[2178] = 12'b000001001110;
		z[2178] = 3'b110;
		y[2179] = 12'b101100110110;
		z[2179] = 3'b100;
		y[2180] = 12'b111110010110;
		z[2180] = 3'b101;
		y[2181] = 12'b110011000011;
		z[2181] = 3'b010;
		y[2182] = 12'b110111100100;
		z[2182] = 3'b100;
		y[2183] = 12'b110000010011;
		z[2183] = 3'b111;
		y[2184] = 12'b100000011111;
		z[2184] = 3'b100;
		y[2185] = 12'b111100111011;
		z[2185] = 3'b010;
		y[2186] = 12'b000111111000;
		z[2186] = 3'b110;
		y[2187] = 12'b001011001101;
		z[2187] = 3'b010;
		y[2188] = 12'b110001100100;
		z[2188] = 3'b011;
		y[2189] = 12'b010000110001;
		z[2189] = 3'b001;
		y[2190] = 12'b100111011010;
		z[2190] = 3'b010;
		y[2191] = 12'b100011101011;
		z[2191] = 3'b110;
		y[2192] = 12'b010000111101;
		z[2192] = 3'b000;
		y[2193] = 12'b111101101101;
		z[2193] = 3'b011;
		y[2194] = 12'b100100101111;
		z[2194] = 3'b010;
		y[2195] = 12'b111111110111;
		z[2195] = 3'b010;
		y[2196] = 12'b010111101001;
		z[2196] = 3'b101;
		y[2197] = 12'b000011010011;
		z[2197] = 3'b011;
		y[2198] = 12'b100010101100;
		z[2198] = 3'b100;
		y[2199] = 12'b111011010001;
		z[2199] = 3'b011;
		y[2200] = 12'b110110000011;
		z[2200] = 3'b110;
		y[2201] = 12'b000101110010;
		z[2201] = 3'b010;
		y[2202] = 12'b100101111111;
		z[2202] = 3'b100;
		y[2203] = 12'b100110110101;
		z[2203] = 3'b011;
		y[2204] = 12'b101111000011;
		z[2204] = 3'b101;
		y[2205] = 12'b110110110000;
		z[2205] = 3'b000;
		y[2206] = 12'b101110101110;
		z[2206] = 3'b111;
		y[2207] = 12'b000100010001;
		z[2207] = 3'b011;
		y[2208] = 12'b111000001100;
		z[2208] = 3'b001;
		y[2209] = 12'b011001011100;
		z[2209] = 3'b110;
		y[2210] = 12'b111001010101;
		z[2210] = 3'b001;
		y[2211] = 12'b100101101001;
		z[2211] = 3'b110;
		y[2212] = 12'b100011001100;
		z[2212] = 3'b010;
		y[2213] = 12'b100010011011;
		z[2213] = 3'b011;
		y[2214] = 12'b110000001011;
		z[2214] = 3'b010;
		y[2215] = 12'b101110010100;
		z[2215] = 3'b011;
		y[2216] = 12'b011001000101;
		z[2216] = 3'b101;
		y[2217] = 12'b111110101010;
		z[2217] = 3'b011;
		y[2218] = 12'b100001000111;
		z[2218] = 3'b000;
		y[2219] = 12'b111110000011;
		z[2219] = 3'b010;
		y[2220] = 12'b111101111110;
		z[2220] = 3'b101;
		y[2221] = 12'b111011010010;
		z[2221] = 3'b111;
		y[2222] = 12'b110000001101;
		z[2222] = 3'b110;
		y[2223] = 12'b111101011000;
		z[2223] = 3'b100;
		y[2224] = 12'b101101010001;
		z[2224] = 3'b010;
		y[2225] = 12'b010010000010;
		z[2225] = 3'b100;
		y[2226] = 12'b111101001111;
		z[2226] = 3'b111;
		y[2227] = 12'b010100001100;
		z[2227] = 3'b101;
		y[2228] = 12'b001000111110;
		z[2228] = 3'b101;
		y[2229] = 12'b101100110111;
		z[2229] = 3'b010;
		y[2230] = 12'b000111011010;
		z[2230] = 3'b001;
		y[2231] = 12'b001101111011;
		z[2231] = 3'b101;
		y[2232] = 12'b010110011110;
		z[2232] = 3'b011;
		y[2233] = 12'b101100110011;
		z[2233] = 3'b011;
		y[2234] = 12'b100110110100;
		z[2234] = 3'b101;
		y[2235] = 12'b000100010001;
		z[2235] = 3'b100;
		y[2236] = 12'b101000110011;
		z[2236] = 3'b100;
		y[2237] = 12'b000100101101;
		z[2237] = 3'b110;
		y[2238] = 12'b101000001010;
		z[2238] = 3'b010;
		y[2239] = 12'b000010011111;
		z[2239] = 3'b010;
		y[2240] = 12'b010101110010;
		z[2240] = 3'b101;
		y[2241] = 12'b101001100111;
		z[2241] = 3'b011;
		y[2242] = 12'b100100001100;
		z[2242] = 3'b111;
		y[2243] = 12'b001110111110;
		z[2243] = 3'b001;
		y[2244] = 12'b101001011000;
		z[2244] = 3'b111;
		y[2245] = 12'b111010100001;
		z[2245] = 3'b101;
		y[2246] = 12'b010100100010;
		z[2246] = 3'b000;
		y[2247] = 12'b001011011101;
		z[2247] = 3'b010;
		y[2248] = 12'b110100010101;
		z[2248] = 3'b101;
		y[2249] = 12'b100001101101;
		z[2249] = 3'b011;
		y[2250] = 12'b101100010001;
		z[2250] = 3'b111;
		y[2251] = 12'b001011110001;
		z[2251] = 3'b100;
		y[2252] = 12'b001001100010;
		z[2252] = 3'b000;
		y[2253] = 12'b001110101001;
		z[2253] = 3'b011;
		y[2254] = 12'b111100000111;
		z[2254] = 3'b001;
		y[2255] = 12'b110111110001;
		z[2255] = 3'b111;
		y[2256] = 12'b000010110111;
		z[2256] = 3'b000;
		y[2257] = 12'b011100000011;
		z[2257] = 3'b100;
		y[2258] = 12'b100001000111;
		z[2258] = 3'b000;
		y[2259] = 12'b010000011101;
		z[2259] = 3'b011;
		y[2260] = 12'b001111111010;
		z[2260] = 3'b011;
		y[2261] = 12'b100000100110;
		z[2261] = 3'b110;
		y[2262] = 12'b000001100011;
		z[2262] = 3'b110;
		y[2263] = 12'b001111011001;
		z[2263] = 3'b001;
		y[2264] = 12'b011110111000;
		z[2264] = 3'b010;
		y[2265] = 12'b011111101011;
		z[2265] = 3'b111;
		y[2266] = 12'b100110111001;
		z[2266] = 3'b111;
		y[2267] = 12'b110000001001;
		z[2267] = 3'b010;
		y[2268] = 12'b001100001101;
		z[2268] = 3'b111;
		y[2269] = 12'b000111100110;
		z[2269] = 3'b101;
		y[2270] = 12'b011010001110;
		z[2270] = 3'b110;
		y[2271] = 12'b010011101011;
		z[2271] = 3'b001;
		y[2272] = 12'b000100100111;
		z[2272] = 3'b001;
		y[2273] = 12'b001100010100;
		z[2273] = 3'b000;
		y[2274] = 12'b110111000100;
		z[2274] = 3'b001;
		y[2275] = 12'b110010011000;
		z[2275] = 3'b110;
		y[2276] = 12'b000011001111;
		z[2276] = 3'b101;
		y[2277] = 12'b000101100010;
		z[2277] = 3'b100;
		y[2278] = 12'b000101110101;
		z[2278] = 3'b111;
		y[2279] = 12'b000110110010;
		z[2279] = 3'b001;
		y[2280] = 12'b011001001101;
		z[2280] = 3'b100;
		y[2281] = 12'b110100011000;
		z[2281] = 3'b001;
		y[2282] = 12'b111110000101;
		z[2282] = 3'b110;
		y[2283] = 12'b011011011010;
		z[2283] = 3'b011;
		y[2284] = 12'b110011110001;
		z[2284] = 3'b010;
		y[2285] = 12'b001001011111;
		z[2285] = 3'b010;
		y[2286] = 12'b101101011001;
		z[2286] = 3'b001;
		y[2287] = 12'b111111100010;
		z[2287] = 3'b100;
		y[2288] = 12'b000000111110;
		z[2288] = 3'b101;
		y[2289] = 12'b110011101010;
		z[2289] = 3'b101;
		y[2290] = 12'b001101110001;
		z[2290] = 3'b000;
		y[2291] = 12'b001100001000;
		z[2291] = 3'b010;
		y[2292] = 12'b111101100001;
		z[2292] = 3'b110;
		y[2293] = 12'b101011000010;
		z[2293] = 3'b101;
		y[2294] = 12'b111000010011;
		z[2294] = 3'b100;
		y[2295] = 12'b110110101010;
		z[2295] = 3'b101;
		y[2296] = 12'b011101111110;
		z[2296] = 3'b001;
		y[2297] = 12'b011111101100;
		z[2297] = 3'b011;
		y[2298] = 12'b001000101110;
		z[2298] = 3'b101;
		y[2299] = 12'b010101010111;
		z[2299] = 3'b000;
		y[2300] = 12'b011110110001;
		z[2300] = 3'b011;
		y[2301] = 12'b110111011010;
		z[2301] = 3'b011;
		y[2302] = 12'b000110110100;
		z[2302] = 3'b010;
		y[2303] = 12'b011111111101;
		z[2303] = 3'b001;
		y[2304] = 12'b100100010111;
		z[2304] = 3'b110;
		y[2305] = 12'b001000100010;
		z[2305] = 3'b011;
		y[2306] = 12'b010111001010;
		z[2306] = 3'b011;
		y[2307] = 12'b110001010110;
		z[2307] = 3'b110;
		y[2308] = 12'b111010010110;
		z[2308] = 3'b001;
		y[2309] = 12'b110111001010;
		z[2309] = 3'b000;
		y[2310] = 12'b100111010010;
		z[2310] = 3'b011;
		y[2311] = 12'b111111010111;
		z[2311] = 3'b101;
		y[2312] = 12'b111111011101;
		z[2312] = 3'b010;
		y[2313] = 12'b000101010100;
		z[2313] = 3'b100;
		y[2314] = 12'b111000010101;
		z[2314] = 3'b001;
		y[2315] = 12'b110010000010;
		z[2315] = 3'b011;
		y[2316] = 12'b010010101010;
		z[2316] = 3'b111;
		y[2317] = 12'b100011000101;
		z[2317] = 3'b101;
		y[2318] = 12'b001101000100;
		z[2318] = 3'b011;
		y[2319] = 12'b010000000000;
		z[2319] = 3'b000;
		y[2320] = 12'b100111011010;
		z[2320] = 3'b100;
		y[2321] = 12'b001101100010;
		z[2321] = 3'b010;
		y[2322] = 12'b110101111011;
		z[2322] = 3'b110;
		y[2323] = 12'b110110000010;
		z[2323] = 3'b111;
		y[2324] = 12'b001111010111;
		z[2324] = 3'b110;
		y[2325] = 12'b001111110101;
		z[2325] = 3'b111;
		y[2326] = 12'b101100100100;
		z[2326] = 3'b110;
		y[2327] = 12'b001001000101;
		z[2327] = 3'b101;
		y[2328] = 12'b010101011000;
		z[2328] = 3'b010;
		y[2329] = 12'b111101100110;
		z[2329] = 3'b010;
		y[2330] = 12'b111000000100;
		z[2330] = 3'b010;
		y[2331] = 12'b100100000010;
		z[2331] = 3'b100;
		y[2332] = 12'b101111111011;
		z[2332] = 3'b000;
		y[2333] = 12'b101001111001;
		z[2333] = 3'b111;
		y[2334] = 12'b011110011001;
		z[2334] = 3'b010;
		y[2335] = 12'b011001000011;
		z[2335] = 3'b101;
		y[2336] = 12'b101110110100;
		z[2336] = 3'b011;
		y[2337] = 12'b011000011011;
		z[2337] = 3'b011;
		y[2338] = 12'b101111010000;
		z[2338] = 3'b110;
		y[2339] = 12'b110100100111;
		z[2339] = 3'b010;
		y[2340] = 12'b011000101111;
		z[2340] = 3'b111;
		y[2341] = 12'b111010110110;
		z[2341] = 3'b011;
		y[2342] = 12'b000011011011;
		z[2342] = 3'b111;
		y[2343] = 12'b010001101001;
		z[2343] = 3'b000;
		y[2344] = 12'b011001011100;
		z[2344] = 3'b111;
		y[2345] = 12'b101001001000;
		z[2345] = 3'b111;
		y[2346] = 12'b111001011110;
		z[2346] = 3'b100;
		y[2347] = 12'b000001111110;
		z[2347] = 3'b100;
		y[2348] = 12'b010011000010;
		z[2348] = 3'b110;
		y[2349] = 12'b100010111011;
		z[2349] = 3'b001;
		y[2350] = 12'b011101110000;
		z[2350] = 3'b100;
		y[2351] = 12'b110001110000;
		z[2351] = 3'b110;
		y[2352] = 12'b100000001111;
		z[2352] = 3'b010;
		y[2353] = 12'b001100110011;
		z[2353] = 3'b100;
		y[2354] = 12'b111111111011;
		z[2354] = 3'b011;
		y[2355] = 12'b100011111011;
		z[2355] = 3'b001;
		y[2356] = 12'b100101100100;
		z[2356] = 3'b111;
		y[2357] = 12'b100010101010;
		z[2357] = 3'b100;
		y[2358] = 12'b011000101000;
		z[2358] = 3'b111;
		y[2359] = 12'b110101111010;
		z[2359] = 3'b000;
		y[2360] = 12'b110110011110;
		z[2360] = 3'b000;
		y[2361] = 12'b001101110111;
		z[2361] = 3'b100;
		y[2362] = 12'b000010110101;
		z[2362] = 3'b111;
		y[2363] = 12'b100100110101;
		z[2363] = 3'b001;
		y[2364] = 12'b110100100000;
		z[2364] = 3'b110;
		y[2365] = 12'b100010111111;
		z[2365] = 3'b100;
		y[2366] = 12'b011010011100;
		z[2366] = 3'b001;
		y[2367] = 12'b100110100000;
		z[2367] = 3'b011;
		y[2368] = 12'b101101110011;
		z[2368] = 3'b110;
		y[2369] = 12'b001000000000;
		z[2369] = 3'b001;
		y[2370] = 12'b100001111101;
		z[2370] = 3'b100;
		y[2371] = 12'b111100111001;
		z[2371] = 3'b110;
		y[2372] = 12'b000110111111;
		z[2372] = 3'b011;
		y[2373] = 12'b111110100110;
		z[2373] = 3'b011;
		y[2374] = 12'b111110010101;
		z[2374] = 3'b100;
		y[2375] = 12'b000010010101;
		z[2375] = 3'b011;
		y[2376] = 12'b011100001011;
		z[2376] = 3'b110;
		y[2377] = 12'b100110011000;
		z[2377] = 3'b100;
		y[2378] = 12'b101101001011;
		z[2378] = 3'b111;
		y[2379] = 12'b010101110011;
		z[2379] = 3'b110;
		y[2380] = 12'b110000101011;
		z[2380] = 3'b001;
		y[2381] = 12'b110011101111;
		z[2381] = 3'b101;
		y[2382] = 12'b110000011100;
		z[2382] = 3'b001;
		y[2383] = 12'b100001000111;
		z[2383] = 3'b101;
		y[2384] = 12'b000000011101;
		z[2384] = 3'b011;
		y[2385] = 12'b000011111100;
		z[2385] = 3'b100;
		y[2386] = 12'b010001110001;
		z[2386] = 3'b101;
		y[2387] = 12'b111001110000;
		z[2387] = 3'b100;
		y[2388] = 12'b111110000010;
		z[2388] = 3'b001;
		y[2389] = 12'b100010011101;
		z[2389] = 3'b001;
		y[2390] = 12'b000000010100;
		z[2390] = 3'b101;
		y[2391] = 12'b000110000100;
		z[2391] = 3'b101;
		y[2392] = 12'b101010101110;
		z[2392] = 3'b010;
		y[2393] = 12'b011011010011;
		z[2393] = 3'b001;
		y[2394] = 12'b110011101100;
		z[2394] = 3'b001;
		y[2395] = 12'b000110000010;
		z[2395] = 3'b000;
		y[2396] = 12'b101111001010;
		z[2396] = 3'b100;
		y[2397] = 12'b000011001110;
		z[2397] = 3'b011;
		y[2398] = 12'b000011010000;
		z[2398] = 3'b000;
		y[2399] = 12'b010001100000;
		z[2399] = 3'b101;
		y[2400] = 12'b011001010001;
		z[2400] = 3'b001;
		y[2401] = 12'b100100010101;
		z[2401] = 3'b101;
		y[2402] = 12'b111111001011;
		z[2402] = 3'b000;
		y[2403] = 12'b001110001110;
		z[2403] = 3'b011;
		y[2404] = 12'b101101001001;
		z[2404] = 3'b101;
		y[2405] = 12'b010110101111;
		z[2405] = 3'b001;
		y[2406] = 12'b011111000101;
		z[2406] = 3'b001;
		y[2407] = 12'b111111111100;
		z[2407] = 3'b000;
		y[2408] = 12'b111100000010;
		z[2408] = 3'b010;
		y[2409] = 12'b101010001110;
		z[2409] = 3'b000;
		y[2410] = 12'b110101010010;
		z[2410] = 3'b000;
		y[2411] = 12'b110001110010;
		z[2411] = 3'b001;
		y[2412] = 12'b011101010100;
		z[2412] = 3'b110;
		y[2413] = 12'b010011010111;
		z[2413] = 3'b101;
		y[2414] = 12'b100010000101;
		z[2414] = 3'b011;
		y[2415] = 12'b110110011011;
		z[2415] = 3'b000;
		y[2416] = 12'b101011000111;
		z[2416] = 3'b110;
		y[2417] = 12'b010101110001;
		z[2417] = 3'b100;
		y[2418] = 12'b001101101111;
		z[2418] = 3'b111;
		y[2419] = 12'b011001101100;
		z[2419] = 3'b011;
		y[2420] = 12'b110000110011;
		z[2420] = 3'b111;
		y[2421] = 12'b110100100000;
		z[2421] = 3'b000;
		y[2422] = 12'b111000110010;
		z[2422] = 3'b001;
		y[2423] = 12'b101001111110;
		z[2423] = 3'b100;
		y[2424] = 12'b000010010100;
		z[2424] = 3'b101;
		y[2425] = 12'b111110100011;
		z[2425] = 3'b000;
		y[2426] = 12'b001000011010;
		z[2426] = 3'b010;
		y[2427] = 12'b001101010011;
		z[2427] = 3'b000;
		y[2428] = 12'b000000111101;
		z[2428] = 3'b000;
		y[2429] = 12'b001110010111;
		z[2429] = 3'b101;
		y[2430] = 12'b100101000110;
		z[2430] = 3'b010;
		y[2431] = 12'b010100101010;
		z[2431] = 3'b001;
		y[2432] = 12'b101110110000;
		z[2432] = 3'b100;
		y[2433] = 12'b011101011101;
		z[2433] = 3'b111;
		y[2434] = 12'b001110111000;
		z[2434] = 3'b110;
		y[2435] = 12'b111101101011;
		z[2435] = 3'b011;
		y[2436] = 12'b000111000011;
		z[2436] = 3'b101;
		y[2437] = 12'b010110111111;
		z[2437] = 3'b110;
		y[2438] = 12'b000000010010;
		z[2438] = 3'b100;
		y[2439] = 12'b001010101100;
		z[2439] = 3'b010;
		y[2440] = 12'b010001000100;
		z[2440] = 3'b111;
		y[2441] = 12'b111001010000;
		z[2441] = 3'b011;
		y[2442] = 12'b010100100100;
		z[2442] = 3'b111;
		y[2443] = 12'b100010101011;
		z[2443] = 3'b000;
		y[2444] = 12'b101010110000;
		z[2444] = 3'b100;
		y[2445] = 12'b000001111000;
		z[2445] = 3'b101;
		y[2446] = 12'b101111100111;
		z[2446] = 3'b000;
		y[2447] = 12'b010011011001;
		z[2447] = 3'b111;
		y[2448] = 12'b010011111111;
		z[2448] = 3'b101;
		y[2449] = 12'b101001100000;
		z[2449] = 3'b011;
		y[2450] = 12'b100100101100;
		z[2450] = 3'b010;
		y[2451] = 12'b001011100100;
		z[2451] = 3'b010;
		y[2452] = 12'b101001000100;
		z[2452] = 3'b100;
		y[2453] = 12'b111100011000;
		z[2453] = 3'b000;
		y[2454] = 12'b001011100111;
		z[2454] = 3'b101;
		y[2455] = 12'b101101011011;
		z[2455] = 3'b000;
		y[2456] = 12'b101110110111;
		z[2456] = 3'b100;
		y[2457] = 12'b011101101100;
		z[2457] = 3'b000;
		y[2458] = 12'b100011010101;
		z[2458] = 3'b001;
		y[2459] = 12'b111010101110;
		z[2459] = 3'b000;
		y[2460] = 12'b011110010011;
		z[2460] = 3'b111;
		y[2461] = 12'b001010101001;
		z[2461] = 3'b001;
		y[2462] = 12'b010011011010;
		z[2462] = 3'b111;
		y[2463] = 12'b011110101110;
		z[2463] = 3'b000;
		y[2464] = 12'b010000011111;
		z[2464] = 3'b010;
		y[2465] = 12'b000000111000;
		z[2465] = 3'b101;
		y[2466] = 12'b110101000011;
		z[2466] = 3'b001;
		y[2467] = 12'b100100001110;
		z[2467] = 3'b010;
		y[2468] = 12'b110001100101;
		z[2468] = 3'b111;
		y[2469] = 12'b010100110100;
		z[2469] = 3'b001;
		y[2470] = 12'b101010011000;
		z[2470] = 3'b111;
		y[2471] = 12'b001101111010;
		z[2471] = 3'b011;
		y[2472] = 12'b010101111110;
		z[2472] = 3'b001;
		y[2473] = 12'b101110011000;
		z[2473] = 3'b100;
		y[2474] = 12'b111110000000;
		z[2474] = 3'b010;
		y[2475] = 12'b001111010010;
		z[2475] = 3'b101;
		y[2476] = 12'b100010011110;
		z[2476] = 3'b100;
		y[2477] = 12'b011000101001;
		z[2477] = 3'b110;
		y[2478] = 12'b111011000000;
		z[2478] = 3'b111;
		y[2479] = 12'b011111000111;
		z[2479] = 3'b101;
		y[2480] = 12'b111101011001;
		z[2480] = 3'b001;
		y[2481] = 12'b101110001110;
		z[2481] = 3'b010;
		y[2482] = 12'b001001011001;
		z[2482] = 3'b110;
		y[2483] = 12'b111011110001;
		z[2483] = 3'b110;
		y[2484] = 12'b111111011101;
		z[2484] = 3'b110;
		y[2485] = 12'b101111111100;
		z[2485] = 3'b101;
		y[2486] = 12'b110000000100;
		z[2486] = 3'b110;
		y[2487] = 12'b010011111011;
		z[2487] = 3'b000;
		y[2488] = 12'b111100010111;
		z[2488] = 3'b011;
		y[2489] = 12'b100010110110;
		z[2489] = 3'b000;
		y[2490] = 12'b101010000010;
		z[2490] = 3'b000;
		y[2491] = 12'b110101111010;
		z[2491] = 3'b100;
		y[2492] = 12'b011000111011;
		z[2492] = 3'b011;
		y[2493] = 12'b110100011010;
		z[2493] = 3'b010;
		y[2494] = 12'b111100011011;
		z[2494] = 3'b110;
		y[2495] = 12'b011001001110;
		z[2495] = 3'b101;
		y[2496] = 12'b011101110100;
		z[2496] = 3'b001;
		y[2497] = 12'b001101110111;
		z[2497] = 3'b101;
		y[2498] = 12'b001010100100;
		z[2498] = 3'b010;
		y[2499] = 12'b010010010101;
		z[2499] = 3'b011;
		y[2500] = 12'b011001110111;
		z[2500] = 3'b011;
		y[2501] = 12'b000000110001;
		z[2501] = 3'b000;
		y[2502] = 12'b010111001011;
		z[2502] = 3'b001;
		y[2503] = 12'b000011011100;
		z[2503] = 3'b101;
		y[2504] = 12'b000010100111;
		z[2504] = 3'b011;
		y[2505] = 12'b001111101011;
		z[2505] = 3'b001;
		y[2506] = 12'b111110011011;
		z[2506] = 3'b111;
		y[2507] = 12'b001010000010;
		z[2507] = 3'b001;
		y[2508] = 12'b100010110100;
		z[2508] = 3'b110;
		y[2509] = 12'b000011110000;
		z[2509] = 3'b110;
		y[2510] = 12'b111011100100;
		z[2510] = 3'b011;
		y[2511] = 12'b100101000111;
		z[2511] = 3'b011;
		y[2512] = 12'b000000000100;
		z[2512] = 3'b010;
		y[2513] = 12'b011001000001;
		z[2513] = 3'b101;
		y[2514] = 12'b011010100111;
		z[2514] = 3'b011;
		y[2515] = 12'b000101001101;
		z[2515] = 3'b011;
		y[2516] = 12'b001110100011;
		z[2516] = 3'b110;
		y[2517] = 12'b111111000100;
		z[2517] = 3'b000;
		y[2518] = 12'b101011001101;
		z[2518] = 3'b111;
		y[2519] = 12'b100100100001;
		z[2519] = 3'b010;
		y[2520] = 12'b110010001011;
		z[2520] = 3'b001;
		y[2521] = 12'b100000101011;
		z[2521] = 3'b000;
		y[2522] = 12'b010101111101;
		z[2522] = 3'b100;
		y[2523] = 12'b111011110001;
		z[2523] = 3'b001;
		y[2524] = 12'b101011001111;
		z[2524] = 3'b111;
		y[2525] = 12'b010001000101;
		z[2525] = 3'b100;
		y[2526] = 12'b110100101111;
		z[2526] = 3'b011;
		y[2527] = 12'b110001001001;
		z[2527] = 3'b000;
		y[2528] = 12'b100101010001;
		z[2528] = 3'b000;
		y[2529] = 12'b100101001000;
		z[2529] = 3'b010;
		y[2530] = 12'b011001000010;
		z[2530] = 3'b011;
		y[2531] = 12'b010110001001;
		z[2531] = 3'b101;
		y[2532] = 12'b011011000101;
		z[2532] = 3'b100;
		y[2533] = 12'b101111000110;
		z[2533] = 3'b000;
		y[2534] = 12'b110010111000;
		z[2534] = 3'b101;
		y[2535] = 12'b010000101100;
		z[2535] = 3'b101;
		y[2536] = 12'b010101001001;
		z[2536] = 3'b011;
		y[2537] = 12'b001011110101;
		z[2537] = 3'b010;
		y[2538] = 12'b100010100011;
		z[2538] = 3'b000;
		y[2539] = 12'b000111000010;
		z[2539] = 3'b010;
		y[2540] = 12'b000111110010;
		z[2540] = 3'b000;
		y[2541] = 12'b011001101011;
		z[2541] = 3'b101;
		y[2542] = 12'b111110001110;
		z[2542] = 3'b011;
		y[2543] = 12'b110101010001;
		z[2543] = 3'b010;
		y[2544] = 12'b010101001100;
		z[2544] = 3'b111;
		y[2545] = 12'b110011010011;
		z[2545] = 3'b101;
		y[2546] = 12'b100110111000;
		z[2546] = 3'b001;
		y[2547] = 12'b010100000100;
		z[2547] = 3'b000;
		y[2548] = 12'b101110111001;
		z[2548] = 3'b010;
		y[2549] = 12'b010101101111;
		z[2549] = 3'b010;
		y[2550] = 12'b011100100001;
		z[2550] = 3'b100;
		y[2551] = 12'b101111010001;
		z[2551] = 3'b111;
		y[2552] = 12'b100111010110;
		z[2552] = 3'b100;
		y[2553] = 12'b001111000001;
		z[2553] = 3'b001;
		y[2554] = 12'b111010000010;
		z[2554] = 3'b000;
		y[2555] = 12'b100101111111;
		z[2555] = 3'b100;
		y[2556] = 12'b111010011011;
		z[2556] = 3'b001;
		y[2557] = 12'b100110010101;
		z[2557] = 3'b001;
		y[2558] = 12'b100001001000;
		z[2558] = 3'b011;
		y[2559] = 12'b110000011011;
		z[2559] = 3'b110;
		y[2560] = 12'b100101000011;
		z[2560] = 3'b011;
		y[2561] = 12'b011111010111;
		z[2561] = 3'b000;
		y[2562] = 12'b011010111100;
		z[2562] = 3'b111;
		y[2563] = 12'b011010101110;
		z[2563] = 3'b000;
		y[2564] = 12'b101000100010;
		z[2564] = 3'b011;
		y[2565] = 12'b001010111000;
		z[2565] = 3'b011;
		y[2566] = 12'b001000010011;
		z[2566] = 3'b100;
		y[2567] = 12'b101110111110;
		z[2567] = 3'b010;
		y[2568] = 12'b111101110101;
		z[2568] = 3'b101;
		y[2569] = 12'b110001010000;
		z[2569] = 3'b111;
		y[2570] = 12'b010001011001;
		z[2570] = 3'b100;
		y[2571] = 12'b110010011110;
		z[2571] = 3'b101;
		y[2572] = 12'b000010111110;
		z[2572] = 3'b011;
		y[2573] = 12'b010100100111;
		z[2573] = 3'b110;
		y[2574] = 12'b100100110000;
		z[2574] = 3'b101;
		y[2575] = 12'b110100001011;
		z[2575] = 3'b110;
		y[2576] = 12'b011011000100;
		z[2576] = 3'b100;
		y[2577] = 12'b010100001000;
		z[2577] = 3'b000;
		y[2578] = 12'b000010010101;
		z[2578] = 3'b010;
		y[2579] = 12'b100111101010;
		z[2579] = 3'b101;
		y[2580] = 12'b101010001001;
		z[2580] = 3'b011;
		y[2581] = 12'b111111010110;
		z[2581] = 3'b101;
		y[2582] = 12'b000001001010;
		z[2582] = 3'b000;
		y[2583] = 12'b011111100001;
		z[2583] = 3'b011;
		y[2584] = 12'b110110101010;
		z[2584] = 3'b111;
		y[2585] = 12'b101110110110;
		z[2585] = 3'b010;
		y[2586] = 12'b010011001101;
		z[2586] = 3'b010;
		y[2587] = 12'b011110100000;
		z[2587] = 3'b001;
		y[2588] = 12'b110001110011;
		z[2588] = 3'b000;
		y[2589] = 12'b011000001001;
		z[2589] = 3'b101;
		y[2590] = 12'b111000000011;
		z[2590] = 3'b110;
		y[2591] = 12'b100001011001;
		z[2591] = 3'b010;
		y[2592] = 12'b000000110011;
		z[2592] = 3'b111;
		y[2593] = 12'b010001100010;
		z[2593] = 3'b111;
		y[2594] = 12'b011101001101;
		z[2594] = 3'b110;
		y[2595] = 12'b100001011001;
		z[2595] = 3'b010;
		y[2596] = 12'b110101101001;
		z[2596] = 3'b111;
		y[2597] = 12'b100101101010;
		z[2597] = 3'b010;
		y[2598] = 12'b000101010111;
		z[2598] = 3'b010;
		y[2599] = 12'b011100110110;
		z[2599] = 3'b010;
		y[2600] = 12'b100100010001;
		z[2600] = 3'b000;
		y[2601] = 12'b111001011100;
		z[2601] = 3'b010;
		y[2602] = 12'b110111010110;
		z[2602] = 3'b001;
		y[2603] = 12'b001000100100;
		z[2603] = 3'b000;
		y[2604] = 12'b111101101011;
		z[2604] = 3'b001;
		y[2605] = 12'b111011000000;
		z[2605] = 3'b000;
		y[2606] = 12'b011100110110;
		z[2606] = 3'b000;
		y[2607] = 12'b010001110011;
		z[2607] = 3'b011;
		y[2608] = 12'b110000111011;
		z[2608] = 3'b010;
		y[2609] = 12'b001110010010;
		z[2609] = 3'b010;
		y[2610] = 12'b001001011110;
		z[2610] = 3'b110;
		y[2611] = 12'b101000110101;
		z[2611] = 3'b001;
		y[2612] = 12'b100111010000;
		z[2612] = 3'b001;
		y[2613] = 12'b101010001001;
		z[2613] = 3'b101;
		y[2614] = 12'b101001100011;
		z[2614] = 3'b111;
		y[2615] = 12'b110000010000;
		z[2615] = 3'b000;
		y[2616] = 12'b011011110000;
		z[2616] = 3'b000;
		y[2617] = 12'b100101110010;
		z[2617] = 3'b111;
		y[2618] = 12'b001001100111;
		z[2618] = 3'b111;
		y[2619] = 12'b100101011001;
		z[2619] = 3'b110;
		y[2620] = 12'b000101111000;
		z[2620] = 3'b001;
		y[2621] = 12'b011110001100;
		z[2621] = 3'b011;
		y[2622] = 12'b010011101110;
		z[2622] = 3'b111;
		y[2623] = 12'b000111111110;
		z[2623] = 3'b110;
		y[2624] = 12'b010100101101;
		z[2624] = 3'b001;
		y[2625] = 12'b001011110000;
		z[2625] = 3'b110;
		y[2626] = 12'b100001101111;
		z[2626] = 3'b111;
		y[2627] = 12'b100000100100;
		z[2627] = 3'b011;
		y[2628] = 12'b001000010011;
		z[2628] = 3'b010;
		y[2629] = 12'b100100000110;
		z[2629] = 3'b001;
		y[2630] = 12'b110110100011;
		z[2630] = 3'b111;
		y[2631] = 12'b001011111001;
		z[2631] = 3'b011;
		y[2632] = 12'b010000100111;
		z[2632] = 3'b001;
		y[2633] = 12'b011010001101;
		z[2633] = 3'b101;
		y[2634] = 12'b101101100110;
		z[2634] = 3'b100;
		y[2635] = 12'b111000010111;
		z[2635] = 3'b001;
		y[2636] = 12'b110100010111;
		z[2636] = 3'b010;
		y[2637] = 12'b011011010110;
		z[2637] = 3'b111;
		y[2638] = 12'b000001110001;
		z[2638] = 3'b101;
		y[2639] = 12'b111111100001;
		z[2639] = 3'b110;
		y[2640] = 12'b001111101011;
		z[2640] = 3'b000;
		y[2641] = 12'b111010011000;
		z[2641] = 3'b011;
		y[2642] = 12'b001100000010;
		z[2642] = 3'b101;
		y[2643] = 12'b101111111011;
		z[2643] = 3'b001;
		y[2644] = 12'b111100000100;
		z[2644] = 3'b110;
		y[2645] = 12'b001000011010;
		z[2645] = 3'b001;
		y[2646] = 12'b111010011111;
		z[2646] = 3'b010;
		y[2647] = 12'b101001100010;
		z[2647] = 3'b110;
		y[2648] = 12'b000001010010;
		z[2648] = 3'b111;
		y[2649] = 12'b001110111010;
		z[2649] = 3'b010;
		y[2650] = 12'b001111100001;
		z[2650] = 3'b100;
		y[2651] = 12'b011011110101;
		z[2651] = 3'b101;
		y[2652] = 12'b110001001110;
		z[2652] = 3'b001;
		y[2653] = 12'b101101100000;
		z[2653] = 3'b110;
		y[2654] = 12'b101000011101;
		z[2654] = 3'b100;
		y[2655] = 12'b101011101000;
		z[2655] = 3'b110;
		y[2656] = 12'b111110111001;
		z[2656] = 3'b001;
		y[2657] = 12'b010000001000;
		z[2657] = 3'b100;
		y[2658] = 12'b010101000110;
		z[2658] = 3'b001;
		y[2659] = 12'b010110001010;
		z[2659] = 3'b111;
		y[2660] = 12'b010001101101;
		z[2660] = 3'b111;
		y[2661] = 12'b011011001001;
		z[2661] = 3'b101;
		y[2662] = 12'b001111110001;
		z[2662] = 3'b000;
		y[2663] = 12'b100011110001;
		z[2663] = 3'b011;
		y[2664] = 12'b011100011000;
		z[2664] = 3'b111;
		y[2665] = 12'b001111001001;
		z[2665] = 3'b110;
		y[2666] = 12'b111011111111;
		z[2666] = 3'b010;
		y[2667] = 12'b000101001000;
		z[2667] = 3'b010;
		y[2668] = 12'b101101011100;
		z[2668] = 3'b110;
		y[2669] = 12'b111110100110;
		z[2669] = 3'b001;
		y[2670] = 12'b111100000111;
		z[2670] = 3'b010;
		y[2671] = 12'b111101011001;
		z[2671] = 3'b101;
		y[2672] = 12'b101111000110;
		z[2672] = 3'b000;
		y[2673] = 12'b011001101100;
		z[2673] = 3'b111;
		y[2674] = 12'b010110011001;
		z[2674] = 3'b111;
		y[2675] = 12'b000111011100;
		z[2675] = 3'b010;
		y[2676] = 12'b111001111010;
		z[2676] = 3'b101;
		y[2677] = 12'b100011011101;
		z[2677] = 3'b011;
		y[2678] = 12'b111011101111;
		z[2678] = 3'b000;
		y[2679] = 12'b101000110000;
		z[2679] = 3'b001;
		y[2680] = 12'b001110101011;
		z[2680] = 3'b101;
		y[2681] = 12'b101111100110;
		z[2681] = 3'b001;
		y[2682] = 12'b011010011111;
		z[2682] = 3'b011;
		y[2683] = 12'b111101100100;
		z[2683] = 3'b111;
		y[2684] = 12'b111000110010;
		z[2684] = 3'b000;
		y[2685] = 12'b000001000111;
		z[2685] = 3'b010;
		y[2686] = 12'b110101101110;
		z[2686] = 3'b110;
		y[2687] = 12'b011011110010;
		z[2687] = 3'b001;
		y[2688] = 12'b110111011010;
		z[2688] = 3'b100;
		y[2689] = 12'b001000110111;
		z[2689] = 3'b100;
		y[2690] = 12'b110100100011;
		z[2690] = 3'b001;
		y[2691] = 12'b101111110101;
		z[2691] = 3'b010;
		y[2692] = 12'b000000110111;
		z[2692] = 3'b001;
		y[2693] = 12'b101111101011;
		z[2693] = 3'b111;
		y[2694] = 12'b110101111000;
		z[2694] = 3'b101;
		y[2695] = 12'b101000111010;
		z[2695] = 3'b010;
		y[2696] = 12'b110110100100;
		z[2696] = 3'b100;
		y[2697] = 12'b110101010011;
		z[2697] = 3'b001;
		y[2698] = 12'b011010100101;
		z[2698] = 3'b101;
		y[2699] = 12'b100100101110;
		z[2699] = 3'b011;
		y[2700] = 12'b111111010001;
		z[2700] = 3'b011;
		y[2701] = 12'b101011100100;
		z[2701] = 3'b100;
		y[2702] = 12'b000011010010;
		z[2702] = 3'b111;
		y[2703] = 12'b101010001011;
		z[2703] = 3'b000;
		y[2704] = 12'b000101100110;
		z[2704] = 3'b100;
		y[2705] = 12'b111011010011;
		z[2705] = 3'b000;
		y[2706] = 12'b011101110101;
		z[2706] = 3'b000;
		y[2707] = 12'b100110111111;
		z[2707] = 3'b101;
		y[2708] = 12'b011111110001;
		z[2708] = 3'b110;
		y[2709] = 12'b000100001111;
		z[2709] = 3'b000;
		y[2710] = 12'b111011101001;
		z[2710] = 3'b011;
		y[2711] = 12'b011001000011;
		z[2711] = 3'b110;
		y[2712] = 12'b010001010101;
		z[2712] = 3'b100;
		y[2713] = 12'b011001001001;
		z[2713] = 3'b010;
		y[2714] = 12'b001010000111;
		z[2714] = 3'b000;
		y[2715] = 12'b001100011000;
		z[2715] = 3'b010;
		y[2716] = 12'b100111010000;
		z[2716] = 3'b001;
		y[2717] = 12'b110010000100;
		z[2717] = 3'b010;
		y[2718] = 12'b101101110000;
		z[2718] = 3'b011;
		y[2719] = 12'b000100011100;
		z[2719] = 3'b001;
		y[2720] = 12'b000010110101;
		z[2720] = 3'b110;
		y[2721] = 12'b111101101010;
		z[2721] = 3'b000;
		y[2722] = 12'b101011011001;
		z[2722] = 3'b110;
		y[2723] = 12'b011100101011;
		z[2723] = 3'b100;
		y[2724] = 12'b000110000011;
		z[2724] = 3'b010;
		y[2725] = 12'b110001100110;
		z[2725] = 3'b011;
		y[2726] = 12'b001001001011;
		z[2726] = 3'b000;
		y[2727] = 12'b101110111001;
		z[2727] = 3'b101;
		y[2728] = 12'b100000001000;
		z[2728] = 3'b111;
		y[2729] = 12'b100010100010;
		z[2729] = 3'b011;
		y[2730] = 12'b001000000111;
		z[2730] = 3'b100;
		y[2731] = 12'b100111001110;
		z[2731] = 3'b111;
		y[2732] = 12'b011011001100;
		z[2732] = 3'b100;
		y[2733] = 12'b111100011110;
		z[2733] = 3'b101;
		y[2734] = 12'b010100001111;
		z[2734] = 3'b100;
		y[2735] = 12'b100001101001;
		z[2735] = 3'b101;
		y[2736] = 12'b110000001000;
		z[2736] = 3'b001;
		y[2737] = 12'b110010111110;
		z[2737] = 3'b000;
		y[2738] = 12'b010111001000;
		z[2738] = 3'b101;
		y[2739] = 12'b010001011011;
		z[2739] = 3'b011;
		y[2740] = 12'b101010001101;
		z[2740] = 3'b001;
		y[2741] = 12'b000101000010;
		z[2741] = 3'b100;
		y[2742] = 12'b010101111000;
		z[2742] = 3'b110;
		y[2743] = 12'b011001010000;
		z[2743] = 3'b111;
		y[2744] = 12'b100010101101;
		z[2744] = 3'b100;
		y[2745] = 12'b011010000111;
		z[2745] = 3'b101;
		y[2746] = 12'b110111001111;
		z[2746] = 3'b000;
		y[2747] = 12'b001110000010;
		z[2747] = 3'b001;
		y[2748] = 12'b010011001010;
		z[2748] = 3'b100;
		y[2749] = 12'b100010110000;
		z[2749] = 3'b010;
		y[2750] = 12'b011101100111;
		z[2750] = 3'b110;
		y[2751] = 12'b111110011010;
		z[2751] = 3'b011;
		y[2752] = 12'b000100001001;
		z[2752] = 3'b011;
		y[2753] = 12'b000010101011;
		z[2753] = 3'b111;
		y[2754] = 12'b000011001011;
		z[2754] = 3'b110;
		y[2755] = 12'b011110011100;
		z[2755] = 3'b100;
		y[2756] = 12'b100011000011;
		z[2756] = 3'b001;
		y[2757] = 12'b100001110010;
		z[2757] = 3'b000;
		y[2758] = 12'b101001000011;
		z[2758] = 3'b100;
		y[2759] = 12'b010010010101;
		z[2759] = 3'b011;
		y[2760] = 12'b010000100101;
		z[2760] = 3'b000;
		y[2761] = 12'b111101100001;
		z[2761] = 3'b001;
		y[2762] = 12'b111011010110;
		z[2762] = 3'b111;
		y[2763] = 12'b101111110000;
		z[2763] = 3'b000;
		y[2764] = 12'b111101000000;
		z[2764] = 3'b100;
		y[2765] = 12'b010111001111;
		z[2765] = 3'b000;
		y[2766] = 12'b101110110000;
		z[2766] = 3'b111;
		y[2767] = 12'b011101100011;
		z[2767] = 3'b111;
		y[2768] = 12'b101011111111;
		z[2768] = 3'b011;
		y[2769] = 12'b001100011000;
		z[2769] = 3'b111;
		y[2770] = 12'b010101100010;
		z[2770] = 3'b110;
		y[2771] = 12'b011000011000;
		z[2771] = 3'b110;
		y[2772] = 12'b111001010111;
		z[2772] = 3'b100;
		y[2773] = 12'b000100111001;
		z[2773] = 3'b010;
		y[2774] = 12'b100000011011;
		z[2774] = 3'b100;
		y[2775] = 12'b101001110100;
		z[2775] = 3'b011;
		y[2776] = 12'b110100110111;
		z[2776] = 3'b000;
		y[2777] = 12'b000101100110;
		z[2777] = 3'b111;
		y[2778] = 12'b000100010101;
		z[2778] = 3'b110;
		y[2779] = 12'b001110010101;
		z[2779] = 3'b001;
		y[2780] = 12'b011101101110;
		z[2780] = 3'b101;
		y[2781] = 12'b101110010011;
		z[2781] = 3'b100;
		y[2782] = 12'b010001000011;
		z[2782] = 3'b010;
		y[2783] = 12'b011100010010;
		z[2783] = 3'b010;
		y[2784] = 12'b011111000110;
		z[2784] = 3'b110;
		y[2785] = 12'b100000000011;
		z[2785] = 3'b111;
		y[2786] = 12'b000110100001;
		z[2786] = 3'b010;
		y[2787] = 12'b100001011001;
		z[2787] = 3'b010;
		y[2788] = 12'b101000010111;
		z[2788] = 3'b110;
		y[2789] = 12'b111001101101;
		z[2789] = 3'b000;
		y[2790] = 12'b010110101001;
		z[2790] = 3'b000;
		y[2791] = 12'b111110101110;
		z[2791] = 3'b100;
		y[2792] = 12'b111110010000;
		z[2792] = 3'b010;
		y[2793] = 12'b010000010011;
		z[2793] = 3'b001;
		y[2794] = 12'b100110011000;
		z[2794] = 3'b000;
		y[2795] = 12'b010110110001;
		z[2795] = 3'b011;
		y[2796] = 12'b101011001110;
		z[2796] = 3'b100;
		y[2797] = 12'b100111111010;
		z[2797] = 3'b001;
		y[2798] = 12'b000001011111;
		z[2798] = 3'b100;
		y[2799] = 12'b111100100101;
		z[2799] = 3'b001;
		y[2800] = 12'b110100110110;
		z[2800] = 3'b110;
		y[2801] = 12'b110000110100;
		z[2801] = 3'b001;
		y[2802] = 12'b101011001001;
		z[2802] = 3'b100;
		y[2803] = 12'b110111111100;
		z[2803] = 3'b011;
		y[2804] = 12'b010111001001;
		z[2804] = 3'b010;
		y[2805] = 12'b100101000111;
		z[2805] = 3'b111;
		y[2806] = 12'b111000001010;
		z[2806] = 3'b000;
		y[2807] = 12'b101110100101;
		z[2807] = 3'b010;
		y[2808] = 12'b010110101000;
		z[2808] = 3'b000;
		y[2809] = 12'b100110110110;
		z[2809] = 3'b100;
		y[2810] = 12'b110001111100;
		z[2810] = 3'b011;
		y[2811] = 12'b111110110001;
		z[2811] = 3'b010;
		y[2812] = 12'b011101000011;
		z[2812] = 3'b000;
		y[2813] = 12'b011011010000;
		z[2813] = 3'b111;
		y[2814] = 12'b100110001111;
		z[2814] = 3'b100;
		y[2815] = 12'b000011110111;
		z[2815] = 3'b011;
		y[2816] = 12'b100110110000;
		z[2816] = 3'b110;
		y[2817] = 12'b010011000111;
		z[2817] = 3'b011;
		y[2818] = 12'b111000110010;
		z[2818] = 3'b001;
		y[2819] = 12'b111100100010;
		z[2819] = 3'b001;
		y[2820] = 12'b111011101011;
		z[2820] = 3'b010;
		y[2821] = 12'b001101100110;
		z[2821] = 3'b001;
		y[2822] = 12'b011110111011;
		z[2822] = 3'b010;
		y[2823] = 12'b011110100110;
		z[2823] = 3'b001;
		y[2824] = 12'b011111011011;
		z[2824] = 3'b001;
		y[2825] = 12'b001111011101;
		z[2825] = 3'b010;
		y[2826] = 12'b101001110010;
		z[2826] = 3'b001;
		y[2827] = 12'b000110101110;
		z[2827] = 3'b111;
		y[2828] = 12'b101101110111;
		z[2828] = 3'b101;
		y[2829] = 12'b011011101000;
		z[2829] = 3'b111;
		y[2830] = 12'b000111010100;
		z[2830] = 3'b011;
		y[2831] = 12'b001111000111;
		z[2831] = 3'b101;
		y[2832] = 12'b100011011010;
		z[2832] = 3'b100;
		y[2833] = 12'b111101110011;
		z[2833] = 3'b101;
		y[2834] = 12'b011000011101;
		z[2834] = 3'b010;
		y[2835] = 12'b110010111011;
		z[2835] = 3'b111;
		y[2836] = 12'b010011010001;
		z[2836] = 3'b010;
		y[2837] = 12'b000010110010;
		z[2837] = 3'b111;
		y[2838] = 12'b001000100100;
		z[2838] = 3'b001;
		y[2839] = 12'b100101101001;
		z[2839] = 3'b111;
		y[2840] = 12'b100111011000;
		z[2840] = 3'b101;
		y[2841] = 12'b110110100010;
		z[2841] = 3'b010;
		y[2842] = 12'b100101010011;
		z[2842] = 3'b010;
		y[2843] = 12'b001110111010;
		z[2843] = 3'b000;
		y[2844] = 12'b001100011011;
		z[2844] = 3'b101;
		y[2845] = 12'b100100011101;
		z[2845] = 3'b111;
		y[2846] = 12'b101100000101;
		z[2846] = 3'b000;
		y[2847] = 12'b111101011001;
		z[2847] = 3'b100;
		y[2848] = 12'b001101001010;
		z[2848] = 3'b100;
		y[2849] = 12'b111011111011;
		z[2849] = 3'b111;
		y[2850] = 12'b101001111001;
		z[2850] = 3'b101;
		y[2851] = 12'b010101111101;
		z[2851] = 3'b010;
		y[2852] = 12'b110100101011;
		z[2852] = 3'b001;
		y[2853] = 12'b010010010010;
		z[2853] = 3'b100;
		y[2854] = 12'b101110000001;
		z[2854] = 3'b101;
		y[2855] = 12'b010001011011;
		z[2855] = 3'b111;
		y[2856] = 12'b101100100010;
		z[2856] = 3'b001;
		y[2857] = 12'b000011110100;
		z[2857] = 3'b000;
		y[2858] = 12'b010101011110;
		z[2858] = 3'b000;
		y[2859] = 12'b110110000000;
		z[2859] = 3'b110;
		y[2860] = 12'b101111010010;
		z[2860] = 3'b010;
		y[2861] = 12'b101011111100;
		z[2861] = 3'b010;
		y[2862] = 12'b101001110011;
		z[2862] = 3'b000;
		y[2863] = 12'b010011010111;
		z[2863] = 3'b010;
		y[2864] = 12'b011101101100;
		z[2864] = 3'b011;
		y[2865] = 12'b010100011110;
		z[2865] = 3'b010;
		y[2866] = 12'b111000100110;
		z[2866] = 3'b101;
		y[2867] = 12'b011010101011;
		z[2867] = 3'b011;
		y[2868] = 12'b100111010100;
		z[2868] = 3'b010;
		y[2869] = 12'b101001001100;
		z[2869] = 3'b000;
		y[2870] = 12'b111101110011;
		z[2870] = 3'b000;
		y[2871] = 12'b111101011010;
		z[2871] = 3'b001;
		y[2872] = 12'b010101000010;
		z[2872] = 3'b001;
		y[2873] = 12'b010110111000;
		z[2873] = 3'b111;
		y[2874] = 12'b110110010100;
		z[2874] = 3'b010;
		y[2875] = 12'b011110100000;
		z[2875] = 3'b001;
		y[2876] = 12'b100000001011;
		z[2876] = 3'b011;
		y[2877] = 12'b001001001000;
		z[2877] = 3'b011;
		y[2878] = 12'b010101110010;
		z[2878] = 3'b100;
		y[2879] = 12'b100100111100;
		z[2879] = 3'b110;
		y[2880] = 12'b011010101001;
		z[2880] = 3'b001;
		y[2881] = 12'b001010010101;
		z[2881] = 3'b110;
		y[2882] = 12'b011001011111;
		z[2882] = 3'b001;
		y[2883] = 12'b110110011111;
		z[2883] = 3'b100;
		y[2884] = 12'b101011101000;
		z[2884] = 3'b110;
		y[2885] = 12'b001010010100;
		z[2885] = 3'b100;
		y[2886] = 12'b011111111010;
		z[2886] = 3'b011;
		y[2887] = 12'b010101000000;
		z[2887] = 3'b100;
		y[2888] = 12'b010011001111;
		z[2888] = 3'b101;
		y[2889] = 12'b000100001100;
		z[2889] = 3'b001;
		y[2890] = 12'b000111000011;
		z[2890] = 3'b011;
		y[2891] = 12'b001010000111;
		z[2891] = 3'b111;
		y[2892] = 12'b011011011011;
		z[2892] = 3'b111;
		y[2893] = 12'b000101011010;
		z[2893] = 3'b010;
		y[2894] = 12'b010111011100;
		z[2894] = 3'b011;
		y[2895] = 12'b101011111001;
		z[2895] = 3'b110;
		y[2896] = 12'b101110011110;
		z[2896] = 3'b110;
		y[2897] = 12'b010111101110;
		z[2897] = 3'b101;
		y[2898] = 12'b010010011100;
		z[2898] = 3'b101;
		y[2899] = 12'b100000110001;
		z[2899] = 3'b010;
		y[2900] = 12'b010000100011;
		z[2900] = 3'b010;
		y[2901] = 12'b010100011101;
		z[2901] = 3'b111;
		y[2902] = 12'b011110001011;
		z[2902] = 3'b110;
		y[2903] = 12'b101011100000;
		z[2903] = 3'b101;
		y[2904] = 12'b100000100101;
		z[2904] = 3'b100;
		y[2905] = 12'b100101101110;
		z[2905] = 3'b111;
		y[2906] = 12'b000000001000;
		z[2906] = 3'b100;
		y[2907] = 12'b011110001010;
		z[2907] = 3'b100;
		y[2908] = 12'b001000111001;
		z[2908] = 3'b010;
		y[2909] = 12'b001000001100;
		z[2909] = 3'b011;
		y[2910] = 12'b101100110011;
		z[2910] = 3'b101;
		y[2911] = 12'b010111101110;
		z[2911] = 3'b000;
		y[2912] = 12'b110100110101;
		z[2912] = 3'b011;
		y[2913] = 12'b111110000100;
		z[2913] = 3'b101;
		y[2914] = 12'b110101010111;
		z[2914] = 3'b000;
		y[2915] = 12'b111111010001;
		z[2915] = 3'b000;
		y[2916] = 12'b000111001000;
		z[2916] = 3'b000;
		y[2917] = 12'b111111010011;
		z[2917] = 3'b101;
		y[2918] = 12'b010011000010;
		z[2918] = 3'b001;
		y[2919] = 12'b100010000010;
		z[2919] = 3'b100;
		y[2920] = 12'b111100111000;
		z[2920] = 3'b010;
		y[2921] = 12'b010001111111;
		z[2921] = 3'b010;
		y[2922] = 12'b010001011010;
		z[2922] = 3'b110;
		y[2923] = 12'b011011001000;
		z[2923] = 3'b000;
		y[2924] = 12'b001100010011;
		z[2924] = 3'b000;
		y[2925] = 12'b011001110100;
		z[2925] = 3'b100;
		y[2926] = 12'b101100100000;
		z[2926] = 3'b101;
		y[2927] = 12'b110011101001;
		z[2927] = 3'b111;
		y[2928] = 12'b100011100011;
		z[2928] = 3'b001;
		y[2929] = 12'b010010010100;
		z[2929] = 3'b001;
		y[2930] = 12'b101001111111;
		z[2930] = 3'b001;
		y[2931] = 12'b110011110100;
		z[2931] = 3'b001;
		y[2932] = 12'b110000001111;
		z[2932] = 3'b100;
		y[2933] = 12'b100000001011;
		z[2933] = 3'b010;
		y[2934] = 12'b101100001001;
		z[2934] = 3'b010;
		y[2935] = 12'b011011010000;
		z[2935] = 3'b110;
		y[2936] = 12'b111110101111;
		z[2936] = 3'b010;
		y[2937] = 12'b101011010010;
		z[2937] = 3'b011;
		y[2938] = 12'b110111010100;
		z[2938] = 3'b100;
		y[2939] = 12'b011110101011;
		z[2939] = 3'b000;
		y[2940] = 12'b011100001100;
		z[2940] = 3'b110;
		y[2941] = 12'b110111111001;
		z[2941] = 3'b001;
		y[2942] = 12'b001111111110;
		z[2942] = 3'b011;
		y[2943] = 12'b001110111011;
		z[2943] = 3'b000;
		y[2944] = 12'b011000110110;
		z[2944] = 3'b000;
		y[2945] = 12'b100101011011;
		z[2945] = 3'b000;
		y[2946] = 12'b110111111000;
		z[2946] = 3'b111;
		y[2947] = 12'b101100101011;
		z[2947] = 3'b111;
		y[2948] = 12'b011001100000;
		z[2948] = 3'b000;
		y[2949] = 12'b101000001000;
		z[2949] = 3'b010;
		y[2950] = 12'b110000000100;
		z[2950] = 3'b010;
		y[2951] = 12'b101000000110;
		z[2951] = 3'b100;
		y[2952] = 12'b010101111111;
		z[2952] = 3'b010;
		y[2953] = 12'b111111010111;
		z[2953] = 3'b100;
		y[2954] = 12'b110101110111;
		z[2954] = 3'b100;
		y[2955] = 12'b101101000001;
		z[2955] = 3'b010;
		y[2956] = 12'b111001110011;
		z[2956] = 3'b010;
		y[2957] = 12'b110001011001;
		z[2957] = 3'b000;
		y[2958] = 12'b000011101001;
		z[2958] = 3'b101;
		y[2959] = 12'b010010000111;
		z[2959] = 3'b011;
		y[2960] = 12'b011010010010;
		z[2960] = 3'b100;
		y[2961] = 12'b011011001001;
		z[2961] = 3'b010;
		y[2962] = 12'b001110010100;
		z[2962] = 3'b101;
		y[2963] = 12'b011010011010;
		z[2963] = 3'b001;
		y[2964] = 12'b100011110000;
		z[2964] = 3'b000;
		y[2965] = 12'b100001010101;
		z[2965] = 3'b111;
		y[2966] = 12'b011001110111;
		z[2966] = 3'b001;
		y[2967] = 12'b011011111000;
		z[2967] = 3'b011;
		y[2968] = 12'b010111001111;
		z[2968] = 3'b100;
		y[2969] = 12'b111110110101;
		z[2969] = 3'b111;
		y[2970] = 12'b001010010011;
		z[2970] = 3'b101;
		y[2971] = 12'b000011111011;
		z[2971] = 3'b001;
		y[2972] = 12'b010111110101;
		z[2972] = 3'b010;
		y[2973] = 12'b000100111100;
		z[2973] = 3'b111;
		y[2974] = 12'b111000011011;
		z[2974] = 3'b110;
		y[2975] = 12'b111100010110;
		z[2975] = 3'b000;
		y[2976] = 12'b111010001101;
		z[2976] = 3'b110;
		y[2977] = 12'b101001111000;
		z[2977] = 3'b101;
		y[2978] = 12'b101011111011;
		z[2978] = 3'b010;
		y[2979] = 12'b101110100111;
		z[2979] = 3'b110;
		y[2980] = 12'b000011101000;
		z[2980] = 3'b000;
		y[2981] = 12'b100101011110;
		z[2981] = 3'b101;
		y[2982] = 12'b100001101101;
		z[2982] = 3'b100;
		y[2983] = 12'b101101000000;
		z[2983] = 3'b100;
		y[2984] = 12'b001000110001;
		z[2984] = 3'b101;
		y[2985] = 12'b001111010101;
		z[2985] = 3'b111;
		y[2986] = 12'b111001010110;
		z[2986] = 3'b011;
		y[2987] = 12'b100011000010;
		z[2987] = 3'b110;
		y[2988] = 12'b101110000001;
		z[2988] = 3'b001;
		y[2989] = 12'b110100101100;
		z[2989] = 3'b011;
		y[2990] = 12'b101111101001;
		z[2990] = 3'b010;
		y[2991] = 12'b001110111110;
		z[2991] = 3'b001;
		y[2992] = 12'b101010001001;
		z[2992] = 3'b110;
		y[2993] = 12'b010100000100;
		z[2993] = 3'b101;
		y[2994] = 12'b101001011101;
		z[2994] = 3'b001;
		y[2995] = 12'b001000000011;
		z[2995] = 3'b010;
		y[2996] = 12'b011011111100;
		z[2996] = 3'b000;
		y[2997] = 12'b110011011111;
		z[2997] = 3'b010;
		y[2998] = 12'b001111000110;
		z[2998] = 3'b001;
		y[2999] = 12'b010110111101;
		z[2999] = 3'b100;
		y[3000] = 12'b110111101001;
		z[3000] = 3'b110;
		y[3001] = 12'b011000000011;
		z[3001] = 3'b101;
		y[3002] = 12'b111101100110;
		z[3002] = 3'b000;
		y[3003] = 12'b010011001000;
		z[3003] = 3'b010;
		y[3004] = 12'b110111011010;
		z[3004] = 3'b110;
		y[3005] = 12'b101101111110;
		z[3005] = 3'b000;
		y[3006] = 12'b101000111110;
		z[3006] = 3'b100;
		y[3007] = 12'b010110100100;
		z[3007] = 3'b101;
		y[3008] = 12'b001101111001;
		z[3008] = 3'b001;
		y[3009] = 12'b010010110100;
		z[3009] = 3'b110;
		y[3010] = 12'b110010000101;
		z[3010] = 3'b110;
		y[3011] = 12'b011010101101;
		z[3011] = 3'b111;
		y[3012] = 12'b110110101010;
		z[3012] = 3'b000;
		y[3013] = 12'b100010011101;
		z[3013] = 3'b110;
		y[3014] = 12'b011110001011;
		z[3014] = 3'b000;
		y[3015] = 12'b111011010000;
		z[3015] = 3'b101;
		y[3016] = 12'b101101010100;
		z[3016] = 3'b110;
		y[3017] = 12'b010101010110;
		z[3017] = 3'b110;
		y[3018] = 12'b100000111010;
		z[3018] = 3'b101;
		y[3019] = 12'b101010001111;
		z[3019] = 3'b100;
		y[3020] = 12'b001101111000;
		z[3020] = 3'b110;
		y[3021] = 12'b010100000011;
		z[3021] = 3'b000;
		y[3022] = 12'b001010010000;
		z[3022] = 3'b110;
		y[3023] = 12'b110010000101;
		z[3023] = 3'b011;
		y[3024] = 12'b010001011101;
		z[3024] = 3'b101;
		y[3025] = 12'b100111100011;
		z[3025] = 3'b011;
		y[3026] = 12'b110110101100;
		z[3026] = 3'b000;
		y[3027] = 12'b011010010010;
		z[3027] = 3'b100;
		y[3028] = 12'b101110110100;
		z[3028] = 3'b111;
		y[3029] = 12'b000001001000;
		z[3029] = 3'b001;
		y[3030] = 12'b011110110101;
		z[3030] = 3'b111;
		y[3031] = 12'b110110011110;
		z[3031] = 3'b000;
		y[3032] = 12'b110110000110;
		z[3032] = 3'b100;
		y[3033] = 12'b100001101101;
		z[3033] = 3'b010;
		y[3034] = 12'b010100100101;
		z[3034] = 3'b000;
		y[3035] = 12'b000001100001;
		z[3035] = 3'b101;
		y[3036] = 12'b110011000100;
		z[3036] = 3'b100;
		y[3037] = 12'b110111011010;
		z[3037] = 3'b101;
		y[3038] = 12'b101100100001;
		z[3038] = 3'b011;
		y[3039] = 12'b001110101110;
		z[3039] = 3'b011;
		y[3040] = 12'b100101010100;
		z[3040] = 3'b111;
		y[3041] = 12'b111100111100;
		z[3041] = 3'b101;
		y[3042] = 12'b000001000110;
		z[3042] = 3'b101;
		y[3043] = 12'b100110111110;
		z[3043] = 3'b010;
		y[3044] = 12'b110010001010;
		z[3044] = 3'b110;
		y[3045] = 12'b101110101011;
		z[3045] = 3'b000;
		y[3046] = 12'b010100111100;
		z[3046] = 3'b010;
		y[3047] = 12'b001010101010;
		z[3047] = 3'b101;
		y[3048] = 12'b110001111000;
		z[3048] = 3'b100;
		y[3049] = 12'b001001010110;
		z[3049] = 3'b111;
		y[3050] = 12'b101011100011;
		z[3050] = 3'b010;
		y[3051] = 12'b100010001100;
		z[3051] = 3'b000;
		y[3052] = 12'b110011100110;
		z[3052] = 3'b100;
		y[3053] = 12'b000000101010;
		z[3053] = 3'b011;
		y[3054] = 12'b100110001010;
		z[3054] = 3'b011;
		y[3055] = 12'b000101000101;
		z[3055] = 3'b100;
		y[3056] = 12'b100001001110;
		z[3056] = 3'b010;
		y[3057] = 12'b101011110101;
		z[3057] = 3'b101;
		y[3058] = 12'b000110010000;
		z[3058] = 3'b000;
		y[3059] = 12'b100010110001;
		z[3059] = 3'b011;
		y[3060] = 12'b001111011001;
		z[3060] = 3'b010;
		y[3061] = 12'b100100101010;
		z[3061] = 3'b101;
		y[3062] = 12'b101010010101;
		z[3062] = 3'b110;
		y[3063] = 12'b011000110110;
		z[3063] = 3'b110;
		y[3064] = 12'b000010111101;
		z[3064] = 3'b110;
		y[3065] = 12'b100100000111;
		z[3065] = 3'b100;
		y[3066] = 12'b100111100011;
		z[3066] = 3'b111;
		y[3067] = 12'b000000011100;
		z[3067] = 3'b110;
		y[3068] = 12'b011111010010;
		z[3068] = 3'b001;
		y[3069] = 12'b110011011101;
		z[3069] = 3'b010;
		y[3070] = 12'b111010110000;
		z[3070] = 3'b010;
		y[3071] = 12'b110000001111;
		z[3071] = 3'b000;
		y[3072] = 12'b010101111000;
		z[3072] = 3'b101;
		y[3073] = 12'b110010001100;
		z[3073] = 3'b001;
		y[3074] = 12'b000011000110;
		z[3074] = 3'b010;
		y[3075] = 12'b111011010010;
		z[3075] = 3'b000;
		y[3076] = 12'b110110101010;
		z[3076] = 3'b010;
		y[3077] = 12'b001101110001;
		z[3077] = 3'b101;
		y[3078] = 12'b011011000010;
		z[3078] = 3'b101;
		y[3079] = 12'b100110001111;
		z[3079] = 3'b111;
		y[3080] = 12'b111111100000;
		z[3080] = 3'b010;
		y[3081] = 12'b011110101111;
		z[3081] = 3'b001;
		y[3082] = 12'b000111011111;
		z[3082] = 3'b110;
		y[3083] = 12'b011011001011;
		z[3083] = 3'b011;
		y[3084] = 12'b011100110010;
		z[3084] = 3'b101;
		y[3085] = 12'b100000110001;
		z[3085] = 3'b111;
		y[3086] = 12'b110100001111;
		z[3086] = 3'b011;
		y[3087] = 12'b110110100011;
		z[3087] = 3'b010;
		y[3088] = 12'b110001011111;
		z[3088] = 3'b001;
		y[3089] = 12'b101000000011;
		z[3089] = 3'b110;
		y[3090] = 12'b100000001011;
		z[3090] = 3'b001;
		y[3091] = 12'b010001000111;
		z[3091] = 3'b111;
		y[3092] = 12'b111101101001;
		z[3092] = 3'b100;
		y[3093] = 12'b010100001000;
		z[3093] = 3'b000;
		y[3094] = 12'b100100010000;
		z[3094] = 3'b100;
		y[3095] = 12'b101110100111;
		z[3095] = 3'b111;
		y[3096] = 12'b001000111001;
		z[3096] = 3'b000;
		y[3097] = 12'b101100111110;
		z[3097] = 3'b111;
		y[3098] = 12'b011001100100;
		z[3098] = 3'b010;
		y[3099] = 12'b011011000000;
		z[3099] = 3'b010;
		y[3100] = 12'b000000001111;
		z[3100] = 3'b010;
		y[3101] = 12'b000100010011;
		z[3101] = 3'b100;
		y[3102] = 12'b111101101100;
		z[3102] = 3'b100;
		y[3103] = 12'b111000101110;
		z[3103] = 3'b100;
		y[3104] = 12'b011110010001;
		z[3104] = 3'b111;
		y[3105] = 12'b110001110111;
		z[3105] = 3'b010;
		y[3106] = 12'b110010000111;
		z[3106] = 3'b111;
		y[3107] = 12'b100101000101;
		z[3107] = 3'b011;
		y[3108] = 12'b000001010101;
		z[3108] = 3'b100;
		y[3109] = 12'b001001001100;
		z[3109] = 3'b110;
		y[3110] = 12'b100000000111;
		z[3110] = 3'b111;
		y[3111] = 12'b011100011111;
		z[3111] = 3'b010;
		y[3112] = 12'b000011010001;
		z[3112] = 3'b101;
		y[3113] = 12'b001100110101;
		z[3113] = 3'b111;
		y[3114] = 12'b001001011101;
		z[3114] = 3'b100;
		y[3115] = 12'b110011001001;
		z[3115] = 3'b001;
		y[3116] = 12'b100100001001;
		z[3116] = 3'b100;
		y[3117] = 12'b010111001011;
		z[3117] = 3'b001;
		y[3118] = 12'b001100010100;
		z[3118] = 3'b011;
		y[3119] = 12'b111101010101;
		z[3119] = 3'b100;
		y[3120] = 12'b110100100101;
		z[3120] = 3'b101;
		y[3121] = 12'b110101111010;
		z[3121] = 3'b110;
		y[3122] = 12'b001001100110;
		z[3122] = 3'b110;
		y[3123] = 12'b011010110100;
		z[3123] = 3'b011;
		y[3124] = 12'b100100011011;
		z[3124] = 3'b001;
		y[3125] = 12'b111011010010;
		z[3125] = 3'b001;
		y[3126] = 12'b100111011001;
		z[3126] = 3'b111;
		y[3127] = 12'b101011101110;
		z[3127] = 3'b011;
		y[3128] = 12'b010100110010;
		z[3128] = 3'b100;
		y[3129] = 12'b010010000100;
		z[3129] = 3'b010;
		y[3130] = 12'b011101101010;
		z[3130] = 3'b101;
		y[3131] = 12'b000011000001;
		z[3131] = 3'b000;
		y[3132] = 12'b100110011100;
		z[3132] = 3'b011;
		y[3133] = 12'b011100001100;
		z[3133] = 3'b000;
		y[3134] = 12'b111000111011;
		z[3134] = 3'b101;
		y[3135] = 12'b111000100001;
		z[3135] = 3'b100;
		y[3136] = 12'b000100111110;
		z[3136] = 3'b111;
		y[3137] = 12'b101110001100;
		z[3137] = 3'b100;
		y[3138] = 12'b111010100111;
		z[3138] = 3'b001;
		y[3139] = 12'b101111001101;
		z[3139] = 3'b100;
		y[3140] = 12'b110010110101;
		z[3140] = 3'b010;
		y[3141] = 12'b010111001100;
		z[3141] = 3'b000;
		y[3142] = 12'b100100001011;
		z[3142] = 3'b110;
		y[3143] = 12'b110110110011;
		z[3143] = 3'b101;
		y[3144] = 12'b001110010000;
		z[3144] = 3'b110;
		y[3145] = 12'b100110000110;
		z[3145] = 3'b000;
		y[3146] = 12'b101000110111;
		z[3146] = 3'b111;
		y[3147] = 12'b011010100011;
		z[3147] = 3'b011;
		y[3148] = 12'b010010010101;
		z[3148] = 3'b100;
		y[3149] = 12'b100110000100;
		z[3149] = 3'b011;
		y[3150] = 12'b111100111011;
		z[3150] = 3'b100;
		y[3151] = 12'b100000001110;
		z[3151] = 3'b011;
		y[3152] = 12'b000010101000;
		z[3152] = 3'b011;
		y[3153] = 12'b110110001000;
		z[3153] = 3'b111;
		y[3154] = 12'b101110001001;
		z[3154] = 3'b010;
		y[3155] = 12'b001101010111;
		z[3155] = 3'b101;
		y[3156] = 12'b001111100011;
		z[3156] = 3'b011;
		y[3157] = 12'b110101111001;
		z[3157] = 3'b001;
		y[3158] = 12'b101100110111;
		z[3158] = 3'b101;
		y[3159] = 12'b001010000011;
		z[3159] = 3'b100;
		y[3160] = 12'b000101110111;
		z[3160] = 3'b110;
		y[3161] = 12'b010010111101;
		z[3161] = 3'b010;
		y[3162] = 12'b001001110110;
		z[3162] = 3'b001;
		y[3163] = 12'b101101011100;
		z[3163] = 3'b101;
		y[3164] = 12'b010000000100;
		z[3164] = 3'b011;
		y[3165] = 12'b110000001000;
		z[3165] = 3'b010;
		y[3166] = 12'b010010010110;
		z[3166] = 3'b001;
		y[3167] = 12'b001100111010;
		z[3167] = 3'b100;
		y[3168] = 12'b110101010001;
		z[3168] = 3'b011;
		y[3169] = 12'b001011010001;
		z[3169] = 3'b011;
		y[3170] = 12'b011110100110;
		z[3170] = 3'b000;
		y[3171] = 12'b010011101101;
		z[3171] = 3'b101;
		y[3172] = 12'b100000111111;
		z[3172] = 3'b001;
		y[3173] = 12'b010100011000;
		z[3173] = 3'b001;
		y[3174] = 12'b100000110000;
		z[3174] = 3'b101;
		y[3175] = 12'b000111010110;
		z[3175] = 3'b011;
		y[3176] = 12'b010101110110;
		z[3176] = 3'b011;
		y[3177] = 12'b110100000110;
		z[3177] = 3'b010;
		y[3178] = 12'b111100010010;
		z[3178] = 3'b001;
		y[3179] = 12'b001001111101;
		z[3179] = 3'b001;
		y[3180] = 12'b010110010011;
		z[3180] = 3'b010;
		y[3181] = 12'b000110001000;
		z[3181] = 3'b001;
		y[3182] = 12'b111111110011;
		z[3182] = 3'b101;
		y[3183] = 12'b111000101110;
		z[3183] = 3'b110;
		y[3184] = 12'b111110010100;
		z[3184] = 3'b110;
		y[3185] = 12'b001011101010;
		z[3185] = 3'b001;
		y[3186] = 12'b011011010101;
		z[3186] = 3'b011;
		y[3187] = 12'b101100001010;
		z[3187] = 3'b101;
		y[3188] = 12'b100010001111;
		z[3188] = 3'b000;
		y[3189] = 12'b011000100010;
		z[3189] = 3'b100;
		y[3190] = 12'b110000010101;
		z[3190] = 3'b111;
		y[3191] = 12'b110100011111;
		z[3191] = 3'b000;
		y[3192] = 12'b111001000010;
		z[3192] = 3'b011;
		y[3193] = 12'b000111011100;
		z[3193] = 3'b100;
		y[3194] = 12'b011110100000;
		z[3194] = 3'b001;
		y[3195] = 12'b010100011110;
		z[3195] = 3'b001;
		y[3196] = 12'b000001010010;
		z[3196] = 3'b010;
		y[3197] = 12'b110110101000;
		z[3197] = 3'b001;
		y[3198] = 12'b001011010001;
		z[3198] = 3'b001;
		y[3199] = 12'b001010110110;
		z[3199] = 3'b001;
		y[3200] = 12'b111110011000;
		z[3200] = 3'b010;
		y[3201] = 12'b011000001101;
		z[3201] = 3'b111;
		y[3202] = 12'b110110101101;
		z[3202] = 3'b100;
		y[3203] = 12'b100000101100;
		z[3203] = 3'b001;
		y[3204] = 12'b111010101000;
		z[3204] = 3'b101;
		y[3205] = 12'b010000101011;
		z[3205] = 3'b111;
		y[3206] = 12'b000110110111;
		z[3206] = 3'b111;
		y[3207] = 12'b101010001100;
		z[3207] = 3'b101;
		y[3208] = 12'b100101001001;
		z[3208] = 3'b000;
		y[3209] = 12'b011000011100;
		z[3209] = 3'b101;
		y[3210] = 12'b110110111001;
		z[3210] = 3'b110;
		y[3211] = 12'b010010100101;
		z[3211] = 3'b011;
		y[3212] = 12'b101000100110;
		z[3212] = 3'b100;
		y[3213] = 12'b011010000110;
		z[3213] = 3'b111;
		y[3214] = 12'b011111000100;
		z[3214] = 3'b011;
		y[3215] = 12'b111111001010;
		z[3215] = 3'b100;
		y[3216] = 12'b001110101101;
		z[3216] = 3'b011;
		y[3217] = 12'b010010110001;
		z[3217] = 3'b110;
		y[3218] = 12'b100100010011;
		z[3218] = 3'b010;
		y[3219] = 12'b111010100111;
		z[3219] = 3'b011;
		y[3220] = 12'b111001010101;
		z[3220] = 3'b111;
		y[3221] = 12'b111000011101;
		z[3221] = 3'b111;
		y[3222] = 12'b001101101100;
		z[3222] = 3'b001;
		y[3223] = 12'b111100101101;
		z[3223] = 3'b101;
		y[3224] = 12'b111110000011;
		z[3224] = 3'b011;
		y[3225] = 12'b001010000011;
		z[3225] = 3'b100;
		y[3226] = 12'b000010100011;
		z[3226] = 3'b001;
		y[3227] = 12'b000001101011;
		z[3227] = 3'b101;
		y[3228] = 12'b000100011000;
		z[3228] = 3'b011;
		y[3229] = 12'b000011101111;
		z[3229] = 3'b101;
		y[3230] = 12'b110000000011;
		z[3230] = 3'b011;
		y[3231] = 12'b010011111110;
		z[3231] = 3'b000;
		y[3232] = 12'b110101001111;
		z[3232] = 3'b011;
		y[3233] = 12'b000011001111;
		z[3233] = 3'b001;
		y[3234] = 12'b001100011110;
		z[3234] = 3'b101;
		y[3235] = 12'b010101111000;
		z[3235] = 3'b110;
		y[3236] = 12'b110101101101;
		z[3236] = 3'b001;
		y[3237] = 12'b011111001100;
		z[3237] = 3'b010;
		y[3238] = 12'b001100101000;
		z[3238] = 3'b101;
		y[3239] = 12'b100100000000;
		z[3239] = 3'b001;
		y[3240] = 12'b011010111111;
		z[3240] = 3'b100;
		y[3241] = 12'b111001011101;
		z[3241] = 3'b001;
		y[3242] = 12'b110001010110;
		z[3242] = 3'b100;
		y[3243] = 12'b100101000000;
		z[3243] = 3'b010;
		y[3244] = 12'b010110001100;
		z[3244] = 3'b110;
		y[3245] = 12'b100000111110;
		z[3245] = 3'b101;
		y[3246] = 12'b000111010101;
		z[3246] = 3'b111;
		y[3247] = 12'b011011011101;
		z[3247] = 3'b001;
		y[3248] = 12'b100110100010;
		z[3248] = 3'b010;
		y[3249] = 12'b111110111011;
		z[3249] = 3'b010;
		y[3250] = 12'b100000011011;
		z[3250] = 3'b101;
		y[3251] = 12'b001010110010;
		z[3251] = 3'b010;
		y[3252] = 12'b101000110110;
		z[3252] = 3'b011;
		y[3253] = 12'b000001110101;
		z[3253] = 3'b000;
		y[3254] = 12'b111110111001;
		z[3254] = 3'b101;
		y[3255] = 12'b101110110111;
		z[3255] = 3'b000;
		y[3256] = 12'b011110111110;
		z[3256] = 3'b100;
		y[3257] = 12'b000110110110;
		z[3257] = 3'b110;
		y[3258] = 12'b111010110100;
		z[3258] = 3'b001;
		y[3259] = 12'b010111011100;
		z[3259] = 3'b110;
		y[3260] = 12'b011000111100;
		z[3260] = 3'b011;
		y[3261] = 12'b000100111110;
		z[3261] = 3'b001;
		y[3262] = 12'b001100101000;
		z[3262] = 3'b000;
		y[3263] = 12'b001111111101;
		z[3263] = 3'b111;
		y[3264] = 12'b110111111100;
		z[3264] = 3'b010;
		y[3265] = 12'b010111010100;
		z[3265] = 3'b011;
		y[3266] = 12'b011011010110;
		z[3266] = 3'b111;
		y[3267] = 12'b100011001011;
		z[3267] = 3'b100;
		y[3268] = 12'b000011001011;
		z[3268] = 3'b110;
		y[3269] = 12'b110110000111;
		z[3269] = 3'b000;
		y[3270] = 12'b010001011001;
		z[3270] = 3'b111;
		y[3271] = 12'b011001101000;
		z[3271] = 3'b111;
		y[3272] = 12'b111111101001;
		z[3272] = 3'b111;
		y[3273] = 12'b101000001101;
		z[3273] = 3'b110;
		y[3274] = 12'b000001100101;
		z[3274] = 3'b000;
		y[3275] = 12'b001001111000;
		z[3275] = 3'b000;
		y[3276] = 12'b111111101001;
		z[3276] = 3'b010;
		y[3277] = 12'b010101000101;
		z[3277] = 3'b110;
		y[3278] = 12'b010110011000;
		z[3278] = 3'b010;
		y[3279] = 12'b010111011100;
		z[3279] = 3'b111;
		y[3280] = 12'b001010000111;
		z[3280] = 3'b001;
		y[3281] = 12'b111010000000;
		z[3281] = 3'b111;
		y[3282] = 12'b001001001001;
		z[3282] = 3'b101;
		y[3283] = 12'b011001011010;
		z[3283] = 3'b100;
		y[3284] = 12'b000010101111;
		z[3284] = 3'b000;
		y[3285] = 12'b110100010011;
		z[3285] = 3'b110;
		y[3286] = 12'b100010001101;
		z[3286] = 3'b101;
		y[3287] = 12'b001110010110;
		z[3287] = 3'b010;
		y[3288] = 12'b110001100101;
		z[3288] = 3'b100;
		y[3289] = 12'b110111000100;
		z[3289] = 3'b101;
		y[3290] = 12'b010000101110;
		z[3290] = 3'b010;
		y[3291] = 12'b000110101011;
		z[3291] = 3'b101;
		y[3292] = 12'b001001000100;
		z[3292] = 3'b111;
		y[3293] = 12'b101100111011;
		z[3293] = 3'b101;
		y[3294] = 12'b000011111101;
		z[3294] = 3'b110;
		y[3295] = 12'b000111001000;
		z[3295] = 3'b010;
		y[3296] = 12'b001101101000;
		z[3296] = 3'b111;
		y[3297] = 12'b101101110000;
		z[3297] = 3'b000;
		y[3298] = 12'b001000110001;
		z[3298] = 3'b000;
		y[3299] = 12'b001100001110;
		z[3299] = 3'b110;
		y[3300] = 12'b100001100011;
		z[3300] = 3'b010;
		y[3301] = 12'b111110100011;
		z[3301] = 3'b000;
		y[3302] = 12'b101100110100;
		z[3302] = 3'b010;
		y[3303] = 12'b001010110010;
		z[3303] = 3'b001;
		y[3304] = 12'b010100001111;
		z[3304] = 3'b011;
		y[3305] = 12'b100010000010;
		z[3305] = 3'b011;
		y[3306] = 12'b011110011111;
		z[3306] = 3'b000;
		y[3307] = 12'b100110100010;
		z[3307] = 3'b000;
		y[3308] = 12'b101000110000;
		z[3308] = 3'b001;
		y[3309] = 12'b000000100010;
		z[3309] = 3'b111;
		y[3310] = 12'b001010010000;
		z[3310] = 3'b011;
		y[3311] = 12'b001011010110;
		z[3311] = 3'b111;
		y[3312] = 12'b010001010001;
		z[3312] = 3'b101;
		y[3313] = 12'b101011110100;
		z[3313] = 3'b110;
		y[3314] = 12'b010110110011;
		z[3314] = 3'b111;
		y[3315] = 12'b100010001001;
		z[3315] = 3'b110;
		y[3316] = 12'b101110000001;
		z[3316] = 3'b100;
		y[3317] = 12'b001100000000;
		z[3317] = 3'b011;
		y[3318] = 12'b111011000111;
		z[3318] = 3'b010;
		y[3319] = 12'b010010000110;
		z[3319] = 3'b010;
		y[3320] = 12'b111101011000;
		z[3320] = 3'b000;
		y[3321] = 12'b111010010001;
		z[3321] = 3'b110;
		y[3322] = 12'b001100011111;
		z[3322] = 3'b110;
		y[3323] = 12'b001010000101;
		z[3323] = 3'b110;
		y[3324] = 12'b111101100110;
		z[3324] = 3'b101;
		y[3325] = 12'b110111010001;
		z[3325] = 3'b010;
		y[3326] = 12'b110101010001;
		z[3326] = 3'b000;
		y[3327] = 12'b101110101011;
		z[3327] = 3'b000;
		y[3328] = 12'b011101000100;
		z[3328] = 3'b100;
		y[3329] = 12'b000111001011;
		z[3329] = 3'b001;
		y[3330] = 12'b011100101100;
		z[3330] = 3'b111;
		y[3331] = 12'b001001100001;
		z[3331] = 3'b111;
		y[3332] = 12'b101111011101;
		z[3332] = 3'b011;
		y[3333] = 12'b011010100001;
		z[3333] = 3'b001;
		y[3334] = 12'b100001101101;
		z[3334] = 3'b101;
		y[3335] = 12'b010100011000;
		z[3335] = 3'b100;
		y[3336] = 12'b001000110001;
		z[3336] = 3'b101;
		y[3337] = 12'b101110110111;
		z[3337] = 3'b100;
		y[3338] = 12'b001001111100;
		z[3338] = 3'b100;
		y[3339] = 12'b101010111010;
		z[3339] = 3'b100;
		y[3340] = 12'b111111110011;
		z[3340] = 3'b001;
		y[3341] = 12'b001001111011;
		z[3341] = 3'b011;
		y[3342] = 12'b011011111101;
		z[3342] = 3'b001;
		y[3343] = 12'b001100101111;
		z[3343] = 3'b100;
		y[3344] = 12'b001100011110;
		z[3344] = 3'b111;
		y[3345] = 12'b010001111011;
		z[3345] = 3'b001;
		y[3346] = 12'b010011100010;
		z[3346] = 3'b110;
		y[3347] = 12'b110000110111;
		z[3347] = 3'b100;
		y[3348] = 12'b000010011101;
		z[3348] = 3'b101;
		y[3349] = 12'b100010011100;
		z[3349] = 3'b000;
		y[3350] = 12'b000010101110;
		z[3350] = 3'b100;
		y[3351] = 12'b111100100110;
		z[3351] = 3'b000;
		y[3352] = 12'b011011000100;
		z[3352] = 3'b010;
		y[3353] = 12'b011111110000;
		z[3353] = 3'b011;
		y[3354] = 12'b011011101101;
		z[3354] = 3'b100;
		y[3355] = 12'b101000100101;
		z[3355] = 3'b011;
		y[3356] = 12'b010010010011;
		z[3356] = 3'b100;
		y[3357] = 12'b010110011110;
		z[3357] = 3'b110;
		y[3358] = 12'b100001001000;
		z[3358] = 3'b100;
		y[3359] = 12'b101101000110;
		z[3359] = 3'b000;
		y[3360] = 12'b100000010101;
		z[3360] = 3'b110;
		y[3361] = 12'b011110010010;
		z[3361] = 3'b100;
		y[3362] = 12'b101000011100;
		z[3362] = 3'b101;
		y[3363] = 12'b011111011111;
		z[3363] = 3'b001;
		y[3364] = 12'b011101001100;
		z[3364] = 3'b010;
		y[3365] = 12'b111001111010;
		z[3365] = 3'b000;
		y[3366] = 12'b001100100101;
		z[3366] = 3'b101;
		y[3367] = 12'b101011010100;
		z[3367] = 3'b101;
		y[3368] = 12'b111000001110;
		z[3368] = 3'b101;
		y[3369] = 12'b100101000011;
		z[3369] = 3'b111;
		y[3370] = 12'b100011010000;
		z[3370] = 3'b000;
		y[3371] = 12'b101011001110;
		z[3371] = 3'b100;
		y[3372] = 12'b011001000010;
		z[3372] = 3'b010;
		y[3373] = 12'b110001011001;
		z[3373] = 3'b111;
		y[3374] = 12'b100011011010;
		z[3374] = 3'b111;
		y[3375] = 12'b100010000100;
		z[3375] = 3'b111;
		y[3376] = 12'b111101100010;
		z[3376] = 3'b101;
		y[3377] = 12'b011010010100;
		z[3377] = 3'b111;
		y[3378] = 12'b010111000000;
		z[3378] = 3'b000;
		y[3379] = 12'b000010001000;
		z[3379] = 3'b000;
		y[3380] = 12'b010100111010;
		z[3380] = 3'b100;
		y[3381] = 12'b111001001110;
		z[3381] = 3'b001;
		y[3382] = 12'b011000110100;
		z[3382] = 3'b000;
		y[3383] = 12'b010101101100;
		z[3383] = 3'b011;
		y[3384] = 12'b100000110101;
		z[3384] = 3'b110;
		y[3385] = 12'b001011000011;
		z[3385] = 3'b000;
		y[3386] = 12'b010100100000;
		z[3386] = 3'b110;
		y[3387] = 12'b010111011110;
		z[3387] = 3'b100;
		y[3388] = 12'b010011000000;
		z[3388] = 3'b010;
		y[3389] = 12'b100100000100;
		z[3389] = 3'b111;
		y[3390] = 12'b101111001100;
		z[3390] = 3'b100;
		y[3391] = 12'b001110000110;
		z[3391] = 3'b000;
		y[3392] = 12'b011000110101;
		z[3392] = 3'b000;
		y[3393] = 12'b101111110001;
		z[3393] = 3'b100;
		y[3394] = 12'b010100110001;
		z[3394] = 3'b100;
		y[3395] = 12'b100110110011;
		z[3395] = 3'b010;
		y[3396] = 12'b101010010001;
		z[3396] = 3'b100;
		y[3397] = 12'b010111001000;
		z[3397] = 3'b000;
		y[3398] = 12'b101011000001;
		z[3398] = 3'b101;
		y[3399] = 12'b000000000111;
		z[3399] = 3'b010;
		y[3400] = 12'b101011011010;
		z[3400] = 3'b000;
		y[3401] = 12'b010001110101;
		z[3401] = 3'b001;
		y[3402] = 12'b100111011001;
		z[3402] = 3'b001;
		y[3403] = 12'b000111010110;
		z[3403] = 3'b000;
		y[3404] = 12'b111011100100;
		z[3404] = 3'b111;
		y[3405] = 12'b100110001100;
		z[3405] = 3'b111;
		y[3406] = 12'b100111000101;
		z[3406] = 3'b101;
		y[3407] = 12'b000000011001;
		z[3407] = 3'b111;
		y[3408] = 12'b000010011001;
		z[3408] = 3'b000;
		y[3409] = 12'b100101100110;
		z[3409] = 3'b110;
		y[3410] = 12'b101101001110;
		z[3410] = 3'b101;
		y[3411] = 12'b100000111001;
		z[3411] = 3'b000;
		y[3412] = 12'b011000110100;
		z[3412] = 3'b000;
		y[3413] = 12'b001001011000;
		z[3413] = 3'b110;
		y[3414] = 12'b000010010100;
		z[3414] = 3'b000;
		y[3415] = 12'b100110001100;
		z[3415] = 3'b010;
		y[3416] = 12'b000110011000;
		z[3416] = 3'b001;
		y[3417] = 12'b010011110100;
		z[3417] = 3'b101;
		y[3418] = 12'b101101101000;
		z[3418] = 3'b101;
		y[3419] = 12'b011001101000;
		z[3419] = 3'b000;
		y[3420] = 12'b110011111011;
		z[3420] = 3'b110;
		y[3421] = 12'b111000101011;
		z[3421] = 3'b001;
		y[3422] = 12'b110100110100;
		z[3422] = 3'b010;
		y[3423] = 12'b001000100001;
		z[3423] = 3'b110;
		y[3424] = 12'b000010011000;
		z[3424] = 3'b110;
		y[3425] = 12'b111100111010;
		z[3425] = 3'b101;
		y[3426] = 12'b010010111000;
		z[3426] = 3'b000;
		y[3427] = 12'b111011001001;
		z[3427] = 3'b010;
		y[3428] = 12'b101011111100;
		z[3428] = 3'b011;
		y[3429] = 12'b001010100010;
		z[3429] = 3'b010;
		y[3430] = 12'b000000010001;
		z[3430] = 3'b110;
		y[3431] = 12'b100010100001;
		z[3431] = 3'b110;
		y[3432] = 12'b110010100101;
		z[3432] = 3'b100;
		y[3433] = 12'b111000100001;
		z[3433] = 3'b011;
		y[3434] = 12'b010001001010;
		z[3434] = 3'b010;
		y[3435] = 12'b110011110111;
		z[3435] = 3'b010;
		y[3436] = 12'b100011000010;
		z[3436] = 3'b111;
		y[3437] = 12'b110101001000;
		z[3437] = 3'b111;
		y[3438] = 12'b101100001110;
		z[3438] = 3'b111;
		y[3439] = 12'b001110111010;
		z[3439] = 3'b000;
		y[3440] = 12'b001000001111;
		z[3440] = 3'b000;
		y[3441] = 12'b000001100010;
		z[3441] = 3'b010;
		y[3442] = 12'b000100101010;
		z[3442] = 3'b100;
		y[3443] = 12'b010001110110;
		z[3443] = 3'b100;
		y[3444] = 12'b101010001101;
		z[3444] = 3'b111;
		y[3445] = 12'b110011000110;
		z[3445] = 3'b000;
		y[3446] = 12'b111000101110;
		z[3446] = 3'b001;
		y[3447] = 12'b000110000100;
		z[3447] = 3'b110;
		y[3448] = 12'b011011100011;
		z[3448] = 3'b111;
		y[3449] = 12'b110100101111;
		z[3449] = 3'b010;
		y[3450] = 12'b011000010000;
		z[3450] = 3'b111;
		y[3451] = 12'b011110110011;
		z[3451] = 3'b011;
		y[3452] = 12'b101011110010;
		z[3452] = 3'b101;
		y[3453] = 12'b011011010010;
		z[3453] = 3'b111;
		y[3454] = 12'b011000001001;
		z[3454] = 3'b010;
		y[3455] = 12'b001101000100;
		z[3455] = 3'b110;
		y[3456] = 12'b000100110001;
		z[3456] = 3'b111;
		y[3457] = 12'b000001011110;
		z[3457] = 3'b101;
		y[3458] = 12'b101100101110;
		z[3458] = 3'b111;
		y[3459] = 12'b011111111110;
		z[3459] = 3'b111;
		y[3460] = 12'b001111110010;
		z[3460] = 3'b110;
		y[3461] = 12'b101111111111;
		z[3461] = 3'b101;
		y[3462] = 12'b000000101110;
		z[3462] = 3'b101;
		y[3463] = 12'b001110001011;
		z[3463] = 3'b111;
		y[3464] = 12'b111001001000;
		z[3464] = 3'b010;
		y[3465] = 12'b000000011100;
		z[3465] = 3'b100;
		y[3466] = 12'b100010111110;
		z[3466] = 3'b110;
		y[3467] = 12'b100001111000;
		z[3467] = 3'b101;
		y[3468] = 12'b000101000110;
		z[3468] = 3'b111;
		y[3469] = 12'b111001100010;
		z[3469] = 3'b101;
		y[3470] = 12'b110110000111;
		z[3470] = 3'b010;
		y[3471] = 12'b011010000101;
		z[3471] = 3'b000;
		y[3472] = 12'b101111110001;
		z[3472] = 3'b100;
		y[3473] = 12'b100101000000;
		z[3473] = 3'b010;
		y[3474] = 12'b101100001101;
		z[3474] = 3'b000;
		y[3475] = 12'b101010100101;
		z[3475] = 3'b000;
		y[3476] = 12'b010001110101;
		z[3476] = 3'b101;
		y[3477] = 12'b100000101110;
		z[3477] = 3'b101;
		y[3478] = 12'b100111001101;
		z[3478] = 3'b011;
		y[3479] = 12'b000010101000;
		z[3479] = 3'b110;
		y[3480] = 12'b011101110001;
		z[3480] = 3'b000;
		y[3481] = 12'b111111001100;
		z[3481] = 3'b101;
		y[3482] = 12'b111000001111;
		z[3482] = 3'b110;
		y[3483] = 12'b100101100001;
		z[3483] = 3'b110;
		y[3484] = 12'b010111000110;
		z[3484] = 3'b110;
		y[3485] = 12'b100111101011;
		z[3485] = 3'b101;
		y[3486] = 12'b000011000111;
		z[3486] = 3'b101;
		y[3487] = 12'b001100010011;
		z[3487] = 3'b101;
		y[3488] = 12'b011110010100;
		z[3488] = 3'b010;
		y[3489] = 12'b100000011000;
		z[3489] = 3'b111;
		y[3490] = 12'b010010010000;
		z[3490] = 3'b000;
		y[3491] = 12'b001110000000;
		z[3491] = 3'b101;
		y[3492] = 12'b011101100101;
		z[3492] = 3'b001;
		y[3493] = 12'b101001111100;
		z[3493] = 3'b011;
		y[3494] = 12'b101001110001;
		z[3494] = 3'b011;
		y[3495] = 12'b011111000010;
		z[3495] = 3'b110;
		y[3496] = 12'b000001010011;
		z[3496] = 3'b000;
		y[3497] = 12'b101100110000;
		z[3497] = 3'b010;
		y[3498] = 12'b100011001000;
		z[3498] = 3'b001;
		y[3499] = 12'b010101100101;
		z[3499] = 3'b000;
		y[3500] = 12'b100000100100;
		z[3500] = 3'b011;
		y[3501] = 12'b101110101111;
		z[3501] = 3'b111;
		y[3502] = 12'b100010001101;
		z[3502] = 3'b001;
		y[3503] = 12'b111011110011;
		z[3503] = 3'b001;
		y[3504] = 12'b001000000011;
		z[3504] = 3'b110;
		y[3505] = 12'b111111101101;
		z[3505] = 3'b001;
		y[3506] = 12'b001111010010;
		z[3506] = 3'b110;
		y[3507] = 12'b111101011011;
		z[3507] = 3'b000;
		y[3508] = 12'b000011000010;
		z[3508] = 3'b100;
		y[3509] = 12'b110010111110;
		z[3509] = 3'b010;
		y[3510] = 12'b111111110001;
		z[3510] = 3'b000;
		y[3511] = 12'b011011110010;
		z[3511] = 3'b100;
		y[3512] = 12'b110001100101;
		z[3512] = 3'b000;
		y[3513] = 12'b110001110100;
		z[3513] = 3'b001;
		y[3514] = 12'b011110101101;
		z[3514] = 3'b100;
		y[3515] = 12'b001100111111;
		z[3515] = 3'b000;
		y[3516] = 12'b101010010110;
		z[3516] = 3'b001;
		y[3517] = 12'b011011110111;
		z[3517] = 3'b111;
		y[3518] = 12'b001101011010;
		z[3518] = 3'b101;
		y[3519] = 12'b110111010101;
		z[3519] = 3'b111;
		y[3520] = 12'b010011111000;
		z[3520] = 3'b110;
		y[3521] = 12'b100110111101;
		z[3521] = 3'b110;
		y[3522] = 12'b111000001101;
		z[3522] = 3'b111;
		y[3523] = 12'b111010011110;
		z[3523] = 3'b101;
		y[3524] = 12'b001110101111;
		z[3524] = 3'b010;
		y[3525] = 12'b111010011010;
		z[3525] = 3'b010;
		y[3526] = 12'b001011000110;
		z[3526] = 3'b001;
		y[3527] = 12'b011010010001;
		z[3527] = 3'b011;
		y[3528] = 12'b000011011100;
		z[3528] = 3'b101;
		y[3529] = 12'b101101101110;
		z[3529] = 3'b000;
		y[3530] = 12'b001000010110;
		z[3530] = 3'b111;
		y[3531] = 12'b100001010111;
		z[3531] = 3'b001;
		y[3532] = 12'b010010000000;
		z[3532] = 3'b011;
		y[3533] = 12'b001111110101;
		z[3533] = 3'b001;
		y[3534] = 12'b010100100010;
		z[3534] = 3'b010;
		y[3535] = 12'b110000001110;
		z[3535] = 3'b100;
		y[3536] = 12'b101011111010;
		z[3536] = 3'b101;
		y[3537] = 12'b001011110110;
		z[3537] = 3'b111;
		y[3538] = 12'b011000110111;
		z[3538] = 3'b101;
		y[3539] = 12'b010101100001;
		z[3539] = 3'b100;
		y[3540] = 12'b111001111101;
		z[3540] = 3'b000;
		y[3541] = 12'b100101000000;
		z[3541] = 3'b101;
		y[3542] = 12'b010111001100;
		z[3542] = 3'b011;
		y[3543] = 12'b000101000010;
		z[3543] = 3'b000;
		y[3544] = 12'b000011111010;
		z[3544] = 3'b110;
		y[3545] = 12'b011100110000;
		z[3545] = 3'b101;
		y[3546] = 12'b110111011110;
		z[3546] = 3'b111;
		y[3547] = 12'b001100111100;
		z[3547] = 3'b100;
		y[3548] = 12'b000101010011;
		z[3548] = 3'b010;
		y[3549] = 12'b010001111100;
		z[3549] = 3'b011;
		y[3550] = 12'b001010001000;
		z[3550] = 3'b100;
		y[3551] = 12'b000100111011;
		z[3551] = 3'b011;
		y[3552] = 12'b001101110000;
		z[3552] = 3'b110;
		y[3553] = 12'b101100010000;
		z[3553] = 3'b100;
		y[3554] = 12'b101001001011;
		z[3554] = 3'b100;
		y[3555] = 12'b100110011100;
		z[3555] = 3'b101;
		y[3556] = 12'b001100100110;
		z[3556] = 3'b001;
		y[3557] = 12'b101000001001;
		z[3557] = 3'b011;
		y[3558] = 12'b010000011111;
		z[3558] = 3'b111;
		y[3559] = 12'b011000101100;
		z[3559] = 3'b010;
		y[3560] = 12'b111110100110;
		z[3560] = 3'b100;
		y[3561] = 12'b100100101111;
		z[3561] = 3'b100;
		y[3562] = 12'b011101100011;
		z[3562] = 3'b110;
		y[3563] = 12'b110010001000;
		z[3563] = 3'b010;
		y[3564] = 12'b000101001100;
		z[3564] = 3'b010;
		y[3565] = 12'b000001000111;
		z[3565] = 3'b100;
		y[3566] = 12'b000010010101;
		z[3566] = 3'b101;
		y[3567] = 12'b101111000111;
		z[3567] = 3'b001;
		y[3568] = 12'b001001001101;
		z[3568] = 3'b100;
		y[3569] = 12'b100110001101;
		z[3569] = 3'b010;
		y[3570] = 12'b111100001100;
		z[3570] = 3'b011;
		y[3571] = 12'b101111101010;
		z[3571] = 3'b000;
		y[3572] = 12'b000100000000;
		z[3572] = 3'b011;
		y[3573] = 12'b111111011011;
		z[3573] = 3'b001;
		y[3574] = 12'b111010110101;
		z[3574] = 3'b001;
		y[3575] = 12'b001110010011;
		z[3575] = 3'b001;
		y[3576] = 12'b110100001001;
		z[3576] = 3'b101;
		y[3577] = 12'b111110001000;
		z[3577] = 3'b011;
		y[3578] = 12'b101110010100;
		z[3578] = 3'b111;
		y[3579] = 12'b000011000011;
		z[3579] = 3'b110;
		y[3580] = 12'b001111101101;
		z[3580] = 3'b101;
		y[3581] = 12'b001000001010;
		z[3581] = 3'b000;
		y[3582] = 12'b011000010001;
		z[3582] = 3'b100;
		y[3583] = 12'b010010011011;
		z[3583] = 3'b001;
		y[3584] = 12'b111001010001;
		z[3584] = 3'b100;
		y[3585] = 12'b011101000100;
		z[3585] = 3'b011;
		y[3586] = 12'b101011110010;
		z[3586] = 3'b010;
		y[3587] = 12'b111111111011;
		z[3587] = 3'b011;
		y[3588] = 12'b011110011001;
		z[3588] = 3'b100;
		y[3589] = 12'b100100110011;
		z[3589] = 3'b110;
		y[3590] = 12'b101111011110;
		z[3590] = 3'b000;
		y[3591] = 12'b100110111011;
		z[3591] = 3'b110;
		y[3592] = 12'b101010000110;
		z[3592] = 3'b111;
		y[3593] = 12'b001111100000;
		z[3593] = 3'b110;
		y[3594] = 12'b011001111111;
		z[3594] = 3'b001;
		y[3595] = 12'b000000010100;
		z[3595] = 3'b101;
		y[3596] = 12'b101011111010;
		z[3596] = 3'b010;
		y[3597] = 12'b101100111001;
		z[3597] = 3'b110;
		y[3598] = 12'b110001011101;
		z[3598] = 3'b000;
		y[3599] = 12'b110101111111;
		z[3599] = 3'b110;
		y[3600] = 12'b011010011010;
		z[3600] = 3'b000;
		y[3601] = 12'b010110110110;
		z[3601] = 3'b001;
		y[3602] = 12'b000110110001;
		z[3602] = 3'b110;
		y[3603] = 12'b001000110111;
		z[3603] = 3'b101;
		y[3604] = 12'b001000010011;
		z[3604] = 3'b100;
		y[3605] = 12'b000111010010;
		z[3605] = 3'b100;
		y[3606] = 12'b001101000011;
		z[3606] = 3'b110;
		y[3607] = 12'b111010011000;
		z[3607] = 3'b101;
		y[3608] = 12'b011100011101;
		z[3608] = 3'b001;
		y[3609] = 12'b101100111011;
		z[3609] = 3'b000;
		y[3610] = 12'b110111010001;
		z[3610] = 3'b110;
		y[3611] = 12'b010011001110;
		z[3611] = 3'b001;
		y[3612] = 12'b100100011001;
		z[3612] = 3'b110;
		y[3613] = 12'b100101100011;
		z[3613] = 3'b000;
		y[3614] = 12'b000011011010;
		z[3614] = 3'b110;
		y[3615] = 12'b101111101110;
		z[3615] = 3'b011;
		y[3616] = 12'b110000011010;
		z[3616] = 3'b010;
		y[3617] = 12'b000111101100;
		z[3617] = 3'b000;
		y[3618] = 12'b011011010010;
		z[3618] = 3'b110;
		y[3619] = 12'b101000100100;
		z[3619] = 3'b111;
		y[3620] = 12'b000001011000;
		z[3620] = 3'b101;
		y[3621] = 12'b010000011010;
		z[3621] = 3'b001;
		y[3622] = 12'b011101001000;
		z[3622] = 3'b101;
		y[3623] = 12'b110001111000;
		z[3623] = 3'b000;
		y[3624] = 12'b111101110011;
		z[3624] = 3'b011;
		y[3625] = 12'b101011101111;
		z[3625] = 3'b100;
		y[3626] = 12'b001111101101;
		z[3626] = 3'b101;
		y[3627] = 12'b100010100000;
		z[3627] = 3'b011;
		y[3628] = 12'b101001110011;
		z[3628] = 3'b100;
		y[3629] = 12'b001001010111;
		z[3629] = 3'b001;
		y[3630] = 12'b100100101000;
		z[3630] = 3'b100;
		y[3631] = 12'b011011101111;
		z[3631] = 3'b111;
		y[3632] = 12'b011111101111;
		z[3632] = 3'b011;
		y[3633] = 12'b010100100100;
		z[3633] = 3'b010;
		y[3634] = 12'b110110101101;
		z[3634] = 3'b111;
		y[3635] = 12'b100100011011;
		z[3635] = 3'b101;
		y[3636] = 12'b111001101111;
		z[3636] = 3'b100;
		y[3637] = 12'b010100110011;
		z[3637] = 3'b100;
		y[3638] = 12'b111011001101;
		z[3638] = 3'b111;
		y[3639] = 12'b110110001001;
		z[3639] = 3'b000;
		y[3640] = 12'b011011111010;
		z[3640] = 3'b111;
		y[3641] = 12'b010011001111;
		z[3641] = 3'b000;
		y[3642] = 12'b100110101011;
		z[3642] = 3'b111;
		y[3643] = 12'b110111110011;
		z[3643] = 3'b111;
		y[3644] = 12'b110111101101;
		z[3644] = 3'b110;
		y[3645] = 12'b110001011110;
		z[3645] = 3'b101;
		y[3646] = 12'b111100101101;
		z[3646] = 3'b000;
		y[3647] = 12'b001111110001;
		z[3647] = 3'b010;
		y[3648] = 12'b111100011101;
		z[3648] = 3'b011;
		y[3649] = 12'b000001001101;
		z[3649] = 3'b101;
		y[3650] = 12'b110010101100;
		z[3650] = 3'b000;
		y[3651] = 12'b101110011101;
		z[3651] = 3'b101;
		y[3652] = 12'b111010010111;
		z[3652] = 3'b111;
		y[3653] = 12'b011110110001;
		z[3653] = 3'b110;
		y[3654] = 12'b100101011111;
		z[3654] = 3'b110;
		y[3655] = 12'b010100000011;
		z[3655] = 3'b111;
		y[3656] = 12'b000010000011;
		z[3656] = 3'b111;
		y[3657] = 12'b000010101010;
		z[3657] = 3'b010;
		y[3658] = 12'b011010011010;
		z[3658] = 3'b100;
		y[3659] = 12'b010110001011;
		z[3659] = 3'b110;
		y[3660] = 12'b010010010000;
		z[3660] = 3'b100;
		y[3661] = 12'b111001110101;
		z[3661] = 3'b110;
		y[3662] = 12'b101110101000;
		z[3662] = 3'b100;
		y[3663] = 12'b011011011110;
		z[3663] = 3'b111;
		y[3664] = 12'b110000111100;
		z[3664] = 3'b000;
		y[3665] = 12'b000011100011;
		z[3665] = 3'b011;
		y[3666] = 12'b001011101111;
		z[3666] = 3'b001;
		y[3667] = 12'b010100010100;
		z[3667] = 3'b010;
		y[3668] = 12'b111010000010;
		z[3668] = 3'b000;
		y[3669] = 12'b000111010111;
		z[3669] = 3'b111;
		y[3670] = 12'b110011100101;
		z[3670] = 3'b100;
		y[3671] = 12'b010100110011;
		z[3671] = 3'b001;
		y[3672] = 12'b100010011011;
		z[3672] = 3'b111;
		y[3673] = 12'b010001000011;
		z[3673] = 3'b100;
		y[3674] = 12'b010100110000;
		z[3674] = 3'b111;
		y[3675] = 12'b011111100011;
		z[3675] = 3'b010;
		y[3676] = 12'b111100011000;
		z[3676] = 3'b100;
		y[3677] = 12'b110011100110;
		z[3677] = 3'b100;
		y[3678] = 12'b010011111100;
		z[3678] = 3'b110;
		y[3679] = 12'b000001010010;
		z[3679] = 3'b111;
		y[3680] = 12'b001111010100;
		z[3680] = 3'b101;
		y[3681] = 12'b110111000101;
		z[3681] = 3'b111;
		y[3682] = 12'b010110011011;
		z[3682] = 3'b011;
		y[3683] = 12'b100010001010;
		z[3683] = 3'b011;
		y[3684] = 12'b000100010110;
		z[3684] = 3'b010;
		y[3685] = 12'b000001100111;
		z[3685] = 3'b101;
		y[3686] = 12'b011101100110;
		z[3686] = 3'b010;
		y[3687] = 12'b010011110001;
		z[3687] = 3'b101;
		y[3688] = 12'b011100000011;
		z[3688] = 3'b010;
		y[3689] = 12'b110011001001;
		z[3689] = 3'b100;
		y[3690] = 12'b100011111111;
		z[3690] = 3'b011;
		y[3691] = 12'b101111000000;
		z[3691] = 3'b100;
		y[3692] = 12'b111011010111;
		z[3692] = 3'b011;
		y[3693] = 12'b001000001010;
		z[3693] = 3'b000;
		y[3694] = 12'b110000100100;
		z[3694] = 3'b101;
		y[3695] = 12'b111101101001;
		z[3695] = 3'b000;
		y[3696] = 12'b010110011001;
		z[3696] = 3'b110;
		y[3697] = 12'b010110010001;
		z[3697] = 3'b011;
		y[3698] = 12'b011001001111;
		z[3698] = 3'b111;
		y[3699] = 12'b111111110110;
		z[3699] = 3'b110;
		y[3700] = 12'b110000110110;
		z[3700] = 3'b111;
		y[3701] = 12'b100110101000;
		z[3701] = 3'b111;
		y[3702] = 12'b100000011100;
		z[3702] = 3'b010;
		y[3703] = 12'b111111101100;
		z[3703] = 3'b101;
		y[3704] = 12'b010011101010;
		z[3704] = 3'b100;
		y[3705] = 12'b100110001000;
		z[3705] = 3'b011;
		y[3706] = 12'b000010011100;
		z[3706] = 3'b001;
		y[3707] = 12'b011110100101;
		z[3707] = 3'b100;
		y[3708] = 12'b110000001011;
		z[3708] = 3'b000;
		y[3709] = 12'b011010110100;
		z[3709] = 3'b011;
		y[3710] = 12'b001001110110;
		z[3710] = 3'b000;
		y[3711] = 12'b110000110101;
		z[3711] = 3'b010;
		y[3712] = 12'b001100000100;
		z[3712] = 3'b101;
		y[3713] = 12'b100101110000;
		z[3713] = 3'b110;
		y[3714] = 12'b111001111100;
		z[3714] = 3'b111;
		y[3715] = 12'b001010010010;
		z[3715] = 3'b001;
		y[3716] = 12'b100011110011;
		z[3716] = 3'b011;
		y[3717] = 12'b101010010110;
		z[3717] = 3'b001;
		y[3718] = 12'b100100100101;
		z[3718] = 3'b011;
		y[3719] = 12'b100001000000;
		z[3719] = 3'b010;
		y[3720] = 12'b101111001000;
		z[3720] = 3'b001;
		y[3721] = 12'b101101100100;
		z[3721] = 3'b101;
		y[3722] = 12'b110001010010;
		z[3722] = 3'b010;
		y[3723] = 12'b110010001001;
		z[3723] = 3'b011;
		y[3724] = 12'b010000010010;
		z[3724] = 3'b001;
		y[3725] = 12'b100100101110;
		z[3725] = 3'b110;
		y[3726] = 12'b110001001000;
		z[3726] = 3'b101;
		y[3727] = 12'b001000001110;
		z[3727] = 3'b001;
		y[3728] = 12'b000011000110;
		z[3728] = 3'b111;
		y[3729] = 12'b100101101001;
		z[3729] = 3'b010;
		y[3730] = 12'b001010111101;
		z[3730] = 3'b000;
		y[3731] = 12'b101110011111;
		z[3731] = 3'b111;
		y[3732] = 12'b111110100101;
		z[3732] = 3'b001;
		y[3733] = 12'b101010011101;
		z[3733] = 3'b101;
		y[3734] = 12'b111100000100;
		z[3734] = 3'b000;
		y[3735] = 12'b000101010110;
		z[3735] = 3'b000;
		y[3736] = 12'b000001001110;
		z[3736] = 3'b001;
		y[3737] = 12'b111100000110;
		z[3737] = 3'b101;
		y[3738] = 12'b010110010010;
		z[3738] = 3'b001;
		y[3739] = 12'b011010001010;
		z[3739] = 3'b011;
		y[3740] = 12'b001100000100;
		z[3740] = 3'b010;
		y[3741] = 12'b000100101111;
		z[3741] = 3'b011;
		y[3742] = 12'b100101011000;
		z[3742] = 3'b101;
		y[3743] = 12'b110000100011;
		z[3743] = 3'b111;
		y[3744] = 12'b101111101111;
		z[3744] = 3'b110;
		y[3745] = 12'b101111100011;
		z[3745] = 3'b011;
		y[3746] = 12'b001010000011;
		z[3746] = 3'b100;
		y[3747] = 12'b000011110011;
		z[3747] = 3'b100;
		y[3748] = 12'b100001010000;
		z[3748] = 3'b101;
		y[3749] = 12'b111100000010;
		z[3749] = 3'b011;
		y[3750] = 12'b001010010011;
		z[3750] = 3'b111;
		y[3751] = 12'b001101001101;
		z[3751] = 3'b001;
		y[3752] = 12'b100101011001;
		z[3752] = 3'b001;
		y[3753] = 12'b011011011011;
		z[3753] = 3'b010;
		y[3754] = 12'b100100000000;
		z[3754] = 3'b000;
		y[3755] = 12'b011010100101;
		z[3755] = 3'b011;
		y[3756] = 12'b011010101111;
		z[3756] = 3'b110;
		y[3757] = 12'b111000010100;
		z[3757] = 3'b100;
		y[3758] = 12'b100101110010;
		z[3758] = 3'b110;
		y[3759] = 12'b111010110000;
		z[3759] = 3'b100;
		y[3760] = 12'b010000110010;
		z[3760] = 3'b000;
		y[3761] = 12'b111000110111;
		z[3761] = 3'b100;
		y[3762] = 12'b000001111100;
		z[3762] = 3'b010;
		y[3763] = 12'b000100001000;
		z[3763] = 3'b000;
		y[3764] = 12'b011100010011;
		z[3764] = 3'b011;
		y[3765] = 12'b111011101111;
		z[3765] = 3'b000;
		y[3766] = 12'b101000111110;
		z[3766] = 3'b010;
		y[3767] = 12'b000010001110;
		z[3767] = 3'b000;
		y[3768] = 12'b011000101101;
		z[3768] = 3'b101;
		y[3769] = 12'b100010000101;
		z[3769] = 3'b011;
		y[3770] = 12'b000001101100;
		z[3770] = 3'b100;
		y[3771] = 12'b111101101011;
		z[3771] = 3'b100;
		y[3772] = 12'b010010001111;
		z[3772] = 3'b010;
		y[3773] = 12'b010100000111;
		z[3773] = 3'b011;
		y[3774] = 12'b100011111000;
		z[3774] = 3'b100;
		y[3775] = 12'b110101100011;
		z[3775] = 3'b110;
		y[3776] = 12'b011011111011;
		z[3776] = 3'b110;
		y[3777] = 12'b010101001101;
		z[3777] = 3'b100;
		y[3778] = 12'b101100110101;
		z[3778] = 3'b001;
		y[3779] = 12'b010101001001;
		z[3779] = 3'b011;
		y[3780] = 12'b010101011011;
		z[3780] = 3'b011;
		y[3781] = 12'b010001001010;
		z[3781] = 3'b010;
		y[3782] = 12'b010110100101;
		z[3782] = 3'b100;
		y[3783] = 12'b011101110010;
		z[3783] = 3'b000;
		y[3784] = 12'b000011000010;
		z[3784] = 3'b111;
		y[3785] = 12'b111000010111;
		z[3785] = 3'b000;
		y[3786] = 12'b100000101010;
		z[3786] = 3'b011;
		y[3787] = 12'b011010111110;
		z[3787] = 3'b100;
		y[3788] = 12'b010011000000;
		z[3788] = 3'b010;
		y[3789] = 12'b010110000011;
		z[3789] = 3'b000;
		y[3790] = 12'b101101011000;
		z[3790] = 3'b110;
		y[3791] = 12'b100111010111;
		z[3791] = 3'b010;
		y[3792] = 12'b101111001101;
		z[3792] = 3'b100;
		y[3793] = 12'b001010111101;
		z[3793] = 3'b111;
		y[3794] = 12'b001001011101;
		z[3794] = 3'b000;
		y[3795] = 12'b010011000111;
		z[3795] = 3'b010;
		y[3796] = 12'b111000101011;
		z[3796] = 3'b100;
		y[3797] = 12'b000010011110;
		z[3797] = 3'b011;
		y[3798] = 12'b100011000100;
		z[3798] = 3'b011;
		y[3799] = 12'b101111011111;
		z[3799] = 3'b110;
		y[3800] = 12'b110001101101;
		z[3800] = 3'b100;
		y[3801] = 12'b110101101001;
		z[3801] = 3'b100;
		y[3802] = 12'b110110010010;
		z[3802] = 3'b000;
		y[3803] = 12'b000101101011;
		z[3803] = 3'b010;
		y[3804] = 12'b000010001010;
		z[3804] = 3'b010;
		y[3805] = 12'b000101000010;
		z[3805] = 3'b011;
		y[3806] = 12'b000101011011;
		z[3806] = 3'b011;
		y[3807] = 12'b011111111110;
		z[3807] = 3'b101;
		y[3808] = 12'b110111001110;
		z[3808] = 3'b010;
		y[3809] = 12'b000010111010;
		z[3809] = 3'b000;
		y[3810] = 12'b010001100100;
		z[3810] = 3'b001;
		y[3811] = 12'b000110101000;
		z[3811] = 3'b111;
		y[3812] = 12'b111001101101;
		z[3812] = 3'b100;
		y[3813] = 12'b010111111001;
		z[3813] = 3'b110;
		y[3814] = 12'b001110111000;
		z[3814] = 3'b001;
		y[3815] = 12'b101110101000;
		z[3815] = 3'b100;
		y[3816] = 12'b001111001111;
		z[3816] = 3'b110;
		y[3817] = 12'b000000111000;
		z[3817] = 3'b011;
		y[3818] = 12'b101101011111;
		z[3818] = 3'b110;
		y[3819] = 12'b101110110000;
		z[3819] = 3'b111;
		y[3820] = 12'b001010101011;
		z[3820] = 3'b001;
		y[3821] = 12'b110001110000;
		z[3821] = 3'b101;
		y[3822] = 12'b011101011101;
		z[3822] = 3'b001;
		y[3823] = 12'b110010000110;
		z[3823] = 3'b111;
		y[3824] = 12'b010011111010;
		z[3824] = 3'b110;
		y[3825] = 12'b011101110110;
		z[3825] = 3'b010;
		y[3826] = 12'b100000001001;
		z[3826] = 3'b111;
		y[3827] = 12'b000111100101;
		z[3827] = 3'b011;
		y[3828] = 12'b101110111010;
		z[3828] = 3'b111;
		y[3829] = 12'b001011111111;
		z[3829] = 3'b101;
		y[3830] = 12'b110011101101;
		z[3830] = 3'b011;
		y[3831] = 12'b001001111100;
		z[3831] = 3'b110;
		y[3832] = 12'b010100111101;
		z[3832] = 3'b000;
		y[3833] = 12'b101000000001;
		z[3833] = 3'b001;
		y[3834] = 12'b111010100011;
		z[3834] = 3'b111;
		y[3835] = 12'b000100001110;
		z[3835] = 3'b111;
		y[3836] = 12'b010110111000;
		z[3836] = 3'b001;
		y[3837] = 12'b101110011000;
		z[3837] = 3'b101;
		y[3838] = 12'b010110000101;
		z[3838] = 3'b011;
		y[3839] = 12'b011101110001;
		z[3839] = 3'b011;
		y[3840] = 12'b000000111101;
		z[3840] = 3'b100;
		y[3841] = 12'b100000101101;
		z[3841] = 3'b000;
		y[3842] = 12'b101101110101;
		z[3842] = 3'b101;
		y[3843] = 12'b110100110010;
		z[3843] = 3'b111;
		y[3844] = 12'b100011011100;
		z[3844] = 3'b010;
		y[3845] = 12'b110010000010;
		z[3845] = 3'b110;
		y[3846] = 12'b001010101100;
		z[3846] = 3'b010;
		y[3847] = 12'b100000011010;
		z[3847] = 3'b100;
		y[3848] = 12'b111101010101;
		z[3848] = 3'b111;
		y[3849] = 12'b100010100101;
		z[3849] = 3'b110;
		y[3850] = 12'b101111010111;
		z[3850] = 3'b100;
		y[3851] = 12'b111101101010;
		z[3851] = 3'b000;
		y[3852] = 12'b010011101100;
		z[3852] = 3'b001;
		y[3853] = 12'b010000101001;
		z[3853] = 3'b001;
		y[3854] = 12'b100100011011;
		z[3854] = 3'b001;
		y[3855] = 12'b100111111100;
		z[3855] = 3'b001;
		y[3856] = 12'b010101000011;
		z[3856] = 3'b101;
		y[3857] = 12'b001000000001;
		z[3857] = 3'b010;
		y[3858] = 12'b010101010110;
		z[3858] = 3'b011;
		y[3859] = 12'b101000001110;
		z[3859] = 3'b111;
		y[3860] = 12'b000011010111;
		z[3860] = 3'b100;
		y[3861] = 12'b101100110011;
		z[3861] = 3'b001;
		y[3862] = 12'b000100101111;
		z[3862] = 3'b100;
		y[3863] = 12'b110101001010;
		z[3863] = 3'b011;
		y[3864] = 12'b101100011010;
		z[3864] = 3'b001;
		y[3865] = 12'b101111110100;
		z[3865] = 3'b011;
		y[3866] = 12'b010110111011;
		z[3866] = 3'b000;
		y[3867] = 12'b101101100001;
		z[3867] = 3'b000;
		y[3868] = 12'b000000101101;
		z[3868] = 3'b011;
		y[3869] = 12'b011010010000;
		z[3869] = 3'b011;
		y[3870] = 12'b100011010101;
		z[3870] = 3'b011;
		y[3871] = 12'b111111111001;
		z[3871] = 3'b010;
		y[3872] = 12'b001011011000;
		z[3872] = 3'b010;
		y[3873] = 12'b111111110010;
		z[3873] = 3'b100;
		y[3874] = 12'b100100100110;
		z[3874] = 3'b111;
		y[3875] = 12'b100111111000;
		z[3875] = 3'b001;
		y[3876] = 12'b110010001111;
		z[3876] = 3'b111;
		y[3877] = 12'b001101001111;
		z[3877] = 3'b001;
		y[3878] = 12'b100011100100;
		z[3878] = 3'b111;
		y[3879] = 12'b100010011001;
		z[3879] = 3'b111;
		y[3880] = 12'b011100000010;
		z[3880] = 3'b111;
		y[3881] = 12'b001011101101;
		z[3881] = 3'b101;
		y[3882] = 12'b101100010000;
		z[3882] = 3'b101;
		y[3883] = 12'b101010010111;
		z[3883] = 3'b111;
		y[3884] = 12'b011101001010;
		z[3884] = 3'b110;
		y[3885] = 12'b011110111001;
		z[3885] = 3'b000;
		y[3886] = 12'b010100110100;
		z[3886] = 3'b000;
		y[3887] = 12'b101100111110;
		z[3887] = 3'b000;
		y[3888] = 12'b101101111100;
		z[3888] = 3'b101;
		y[3889] = 12'b000100100010;
		z[3889] = 3'b100;
		y[3890] = 12'b011010001100;
		z[3890] = 3'b000;
		y[3891] = 12'b000110110001;
		z[3891] = 3'b111;
		y[3892] = 12'b000111101011;
		z[3892] = 3'b101;
		y[3893] = 12'b000000100011;
		z[3893] = 3'b010;
		y[3894] = 12'b100101100000;
		z[3894] = 3'b100;
		y[3895] = 12'b111100100101;
		z[3895] = 3'b110;
		y[3896] = 12'b110110011001;
		z[3896] = 3'b101;
		y[3897] = 12'b001100100000;
		z[3897] = 3'b011;
		y[3898] = 12'b001011000101;
		z[3898] = 3'b111;
		y[3899] = 12'b110001110000;
		z[3899] = 3'b111;
		y[3900] = 12'b001110000001;
		z[3900] = 3'b111;
		y[3901] = 12'b000111101101;
		z[3901] = 3'b101;
		y[3902] = 12'b110011001000;
		z[3902] = 3'b011;
		y[3903] = 12'b001010111010;
		z[3903] = 3'b001;
		y[3904] = 12'b111000111001;
		z[3904] = 3'b100;
		y[3905] = 12'b010110011000;
		z[3905] = 3'b010;
		y[3906] = 12'b001111010110;
		z[3906] = 3'b010;
		y[3907] = 12'b010000001010;
		z[3907] = 3'b101;
		y[3908] = 12'b010000110110;
		z[3908] = 3'b110;
		y[3909] = 12'b110110100010;
		z[3909] = 3'b100;
		y[3910] = 12'b000110011000;
		z[3910] = 3'b011;
		y[3911] = 12'b011011110011;
		z[3911] = 3'b101;
		y[3912] = 12'b000010101100;
		z[3912] = 3'b100;
		y[3913] = 12'b010000000110;
		z[3913] = 3'b011;
		y[3914] = 12'b011011110110;
		z[3914] = 3'b101;
		y[3915] = 12'b101100111111;
		z[3915] = 3'b110;
		y[3916] = 12'b100110101101;
		z[3916] = 3'b101;
		y[3917] = 12'b100101101001;
		z[3917] = 3'b110;
		y[3918] = 12'b010111111110;
		z[3918] = 3'b100;
		y[3919] = 12'b100001010111;
		z[3919] = 3'b100;
		y[3920] = 12'b011101011101;
		z[3920] = 3'b001;
		y[3921] = 12'b000010111011;
		z[3921] = 3'b110;
		y[3922] = 12'b011001111001;
		z[3922] = 3'b110;
		y[3923] = 12'b010101010010;
		z[3923] = 3'b010;
		y[3924] = 12'b100111000101;
		z[3924] = 3'b000;
		y[3925] = 12'b100110101100;
		z[3925] = 3'b000;
		y[3926] = 12'b001001001110;
		z[3926] = 3'b010;
		y[3927] = 12'b001110000111;
		z[3927] = 3'b000;
		y[3928] = 12'b001110101100;
		z[3928] = 3'b010;
		y[3929] = 12'b100000001000;
		z[3929] = 3'b011;
		y[3930] = 12'b110011011100;
		z[3930] = 3'b110;
		y[3931] = 12'b000000110111;
		z[3931] = 3'b101;
		y[3932] = 12'b000110001011;
		z[3932] = 3'b001;
		y[3933] = 12'b100100111101;
		z[3933] = 3'b011;
		y[3934] = 12'b111010100111;
		z[3934] = 3'b001;
		y[3935] = 12'b100011100000;
		z[3935] = 3'b001;
		y[3936] = 12'b011001110111;
		z[3936] = 3'b011;
		y[3937] = 12'b000010111110;
		z[3937] = 3'b110;
		y[3938] = 12'b101011100001;
		z[3938] = 3'b011;
		y[3939] = 12'b100000011111;
		z[3939] = 3'b001;
		y[3940] = 12'b010011101001;
		z[3940] = 3'b100;
		y[3941] = 12'b101101111001;
		z[3941] = 3'b101;
		y[3942] = 12'b100011110000;
		z[3942] = 3'b111;
		y[3943] = 12'b110001100010;
		z[3943] = 3'b110;
		y[3944] = 12'b100000101001;
		z[3944] = 3'b100;
		y[3945] = 12'b000001110111;
		z[3945] = 3'b011;
		y[3946] = 12'b100011011000;
		z[3946] = 3'b101;
		y[3947] = 12'b101010100010;
		z[3947] = 3'b011;
		y[3948] = 12'b100001001100;
		z[3948] = 3'b010;
		y[3949] = 12'b001001101101;
		z[3949] = 3'b101;
		y[3950] = 12'b010101110100;
		z[3950] = 3'b101;
		y[3951] = 12'b111100011010;
		z[3951] = 3'b111;
		y[3952] = 12'b000100000101;
		z[3952] = 3'b001;
		y[3953] = 12'b011100001100;
		z[3953] = 3'b100;
		y[3954] = 12'b111111101001;
		z[3954] = 3'b000;
		y[3955] = 12'b100101111101;
		z[3955] = 3'b110;
		y[3956] = 12'b010111011011;
		z[3956] = 3'b101;
		y[3957] = 12'b100000111000;
		z[3957] = 3'b111;
		y[3958] = 12'b010001110000;
		z[3958] = 3'b100;
		y[3959] = 12'b101001000111;
		z[3959] = 3'b100;
		y[3960] = 12'b101000101100;
		z[3960] = 3'b101;
		y[3961] = 12'b011101010000;
		z[3961] = 3'b111;
		y[3962] = 12'b110001010100;
		z[3962] = 3'b011;
		y[3963] = 12'b000001011101;
		z[3963] = 3'b011;
		y[3964] = 12'b110111110011;
		z[3964] = 3'b101;
		y[3965] = 12'b110100010001;
		z[3965] = 3'b001;
		y[3966] = 12'b001011101000;
		z[3966] = 3'b101;
		y[3967] = 12'b011100100001;
		z[3967] = 3'b001;
		y[3968] = 12'b100000110111;
		z[3968] = 3'b010;
		y[3969] = 12'b011001001110;
		z[3969] = 3'b010;
		y[3970] = 12'b100010101011;
		z[3970] = 3'b010;
		y[3971] = 12'b011111000110;
		z[3971] = 3'b100;
		y[3972] = 12'b110100110010;
		z[3972] = 3'b101;
		y[3973] = 12'b000010001000;
		z[3973] = 3'b010;
		y[3974] = 12'b001000111000;
		z[3974] = 3'b010;
		y[3975] = 12'b110111111001;
		z[3975] = 3'b111;
		y[3976] = 12'b110011110010;
		z[3976] = 3'b011;
		y[3977] = 12'b101011001111;
		z[3977] = 3'b110;
		y[3978] = 12'b011100101000;
		z[3978] = 3'b100;
		y[3979] = 12'b011110111100;
		z[3979] = 3'b110;
		y[3980] = 12'b000000101100;
		z[3980] = 3'b000;
		y[3981] = 12'b100110001100;
		z[3981] = 3'b000;
		y[3982] = 12'b011001010000;
		z[3982] = 3'b110;
		y[3983] = 12'b000101001001;
		z[3983] = 3'b100;
		y[3984] = 12'b100001011111;
		z[3984] = 3'b111;
		y[3985] = 12'b010011111000;
		z[3985] = 3'b110;
		y[3986] = 12'b111010111100;
		z[3986] = 3'b001;
		y[3987] = 12'b000111101100;
		z[3987] = 3'b101;
		y[3988] = 12'b110001000110;
		z[3988] = 3'b011;
		y[3989] = 12'b101100000000;
		z[3989] = 3'b110;
		y[3990] = 12'b100111000110;
		z[3990] = 3'b100;
		y[3991] = 12'b000101110110;
		z[3991] = 3'b111;
		y[3992] = 12'b101011110000;
		z[3992] = 3'b000;
		y[3993] = 12'b100010100000;
		z[3993] = 3'b100;
		y[3994] = 12'b100001111110;
		z[3994] = 3'b010;
		y[3995] = 12'b010001100011;
		z[3995] = 3'b011;
		y[3996] = 12'b010001110001;
		z[3996] = 3'b110;
		y[3997] = 12'b000000101011;
		z[3997] = 3'b110;
		y[3998] = 12'b010110000000;
		z[3998] = 3'b011;
		y[3999] = 12'b000100100010;
		z[3999] = 3'b110;
	
		//initialize stimulus_list with zeros
        y_list = 0;
        z_list = 0;
        
        //concatenate all stimulus generated above 
        for(i = 0; i < `STIMULUS_WIDTH; i = i + 1) begin
            y_list = y_list + y[i];
            z_list = z_list + z[i];
            if(i < (`STIMULUS_WIDTH - 1)) begin
                y_list = y_list << `DATA_WIDTH;
                z_list = z_list << `CTRL_WIDTH;
            end 
            //$write("y_list = %b \n", y_list);
            //$write("z_list = %b \n", z_list);
        end
	end
endmodule
