module test;
    
tester tester();

endmodule

