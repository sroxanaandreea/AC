module fsm_trecere(
    output reg p_rosu,      // red for pedestrians
    output reg p_verde,     // green for pedestrians
    output reg m_rosu,      // red for cars
    output reg m_galben,    // yellow for cars
    output reg m_verde,     // green for cars
    output reg [7:0] T,     // timeout count
    input done,             // timeout expired
    input clk);             // clock input

// TODO: Implementarea trecerii de pietoni semaforizata

endmodule