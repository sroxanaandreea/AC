`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:16:24 10/19/2020 
// Design Name: 
// Module Name:    demux1_4 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module demux1_4(
    input in,
    input [1:0] sel,
    output out1,
    output out2,
    output out3,
    output out4
    );

//TODO implementarea functionalitatii unui demultiplexor

endmodule
