module adder6(output[6:0] sum,input[5:0]a,b);

assign sum a + b;
endmodule
