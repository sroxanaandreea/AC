module trecere(
    output p_rosu,          // red for pedestrians
    output p_verde,         // green for pedestrians
    output m_rosu,          // red for cars
    output m_galben,        // yellow for cars
    output m_verde,         // green for cars
    input clk);             // clock input

// TODO: Realizati conexiunile cu automatul de stari

endmodule
